-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
package iu_exec_global_package is -- 
  constant ACCESS_ASR : std_logic_vector(2 downto 0) := "101";
  constant ACCESS_PSR : std_logic_vector(2 downto 0) := "001";
  constant ACCESS_REG : std_logic_vector(2 downto 0) := "110";
  constant ACCESS_TBR : std_logic_vector(2 downto 0) := "010";
  constant ACCESS_WIM : std_logic_vector(2 downto 0) := "011";
  constant ACCESS_Y : std_logic_vector(2 downto 0) := "100";
  constant ALU_INSTR : std_logic_vector(2 downto 0) := "010";
  constant ANNUL_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000000000000001000";
  constant ANNUL_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000000011";
  constant ASI_AJIT_BRIDGE_CONFIG : std_logic_vector(7 downto 0) := "00110000";
  constant ASI_BLOCK_COPY : std_logic_vector(7 downto 0) := "00010111";
  constant ASI_BLOCK_FILL : std_logic_vector(7 downto 0) := "00011111";
  constant ASI_CACHE_DATA_I : std_logic_vector(7 downto 0) := "00001101";
  constant ASI_CACHE_DATA_I_D : std_logic_vector(7 downto 0) := "00001111";
  constant ASI_CACHE_TAG_I : std_logic_vector(7 downto 0) := "00001100";
  constant ASI_CACHE_TAG_I_D : std_logic_vector(7 downto 0) := "00001110";
  constant ASI_FLUSH_I_CONTEXT : std_logic_vector(7 downto 0) := "00011011";
  constant ASI_FLUSH_I_D_CONTEXT : std_logic_vector(7 downto 0) := "00010011";
  constant ASI_FLUSH_I_D_PAGE : std_logic_vector(7 downto 0) := "00010000";
  constant ASI_FLUSH_I_D_REGION : std_logic_vector(7 downto 0) := "00010010";
  constant ASI_FLUSH_I_D_SEGMENT : std_logic_vector(7 downto 0) := "00010001";
  constant ASI_FLUSH_I_D_USER : std_logic_vector(7 downto 0) := "00010100";
  constant ASI_FLUSH_I_PAGE : std_logic_vector(7 downto 0) := "00011000";
  constant ASI_FLUSH_I_REGION : std_logic_vector(7 downto 0) := "00011010";
  constant ASI_FLUSH_I_SEGMENT : std_logic_vector(7 downto 0) := "00011001";
  constant ASI_FLUSH_I_USER : std_logic_vector(7 downto 0) := "00011100";
  constant ASI_MMU_DIAGNOSTIC_I : std_logic_vector(7 downto 0) := "00000101";
  constant ASI_MMU_DIAGNOSTIC_IO : std_logic_vector(7 downto 0) := "00000111";
  constant ASI_MMU_DIAGNOSTIC_I_D : std_logic_vector(7 downto 0) := "00000110";
  constant ASI_MMU_FLUSH_PROBE : std_logic_vector(7 downto 0) := "00000011";
  constant ASI_MMU_REGISTER : std_logic_vector(7 downto 0) := "00000100";
  constant ASI_SUPERVISOR_DATA : std_logic_vector(7 downto 0) := "00001011";
  constant ASI_SUPERVISOR_INSTRUCTION : std_logic_vector(7 downto 0) := "00001001";
  constant ASI_USER_DATA : std_logic_vector(7 downto 0) := "00001010";
  constant ASI_USER_INSTRUCTION : std_logic_vector(7 downto 0) := "00001000";
  constant BLOCK_READ : std_logic_vector(0 downto 0) := "1";
  constant CACHE_ARRAY_NOP : std_logic_vector(2 downto 0) := "011";
  constant CACHE_ARRAY_PASS_THROUGH : std_logic_vector(2 downto 0) := "100";
  constant CACHE_ARRAY_READ_DWORD : std_logic_vector(2 downto 0) := "001";
  constant CACHE_ARRAY_WRITE_DWORD : std_logic_vector(2 downto 0) := "010";
  constant CACHE_TAG_CLEAR_ALL : std_logic_vector(2 downto 0) := "100";
  constant CACHE_TAG_CLEAR_LINE : std_logic_vector(2 downto 0) := "011";
  constant CACHE_TAG_INSERT : std_logic_vector(2 downto 0) := "010";
  constant CACHE_TAG_LOOKUP : std_logic_vector(2 downto 0) := "001";
  constant CACHE_TAG_NOP : std_logic_vector(2 downto 0) := "101";
  constant CCU_DBG_BP_HIT : std_logic_vector(7 downto 0) := "00000010";
  constant CCU_DBG_CONNECT_RQST : std_logic_vector(7 downto 0) := "00000001";
  constant CCU_DBG_ERROR : std_logic_vector(7 downto 0) := "00000111";
  constant CCU_DBG_ERROR_MODE : std_logic_vector(7 downto 0) := "00000110";
  constant CCU_DBG_OK : std_logic_vector(7 downto 0) := "00001000";
  constant CCU_DBG_READ_RESPONSE : std_logic_vector(7 downto 0) := "00001001";
  constant CCU_DBG_READ_WP_HIT : std_logic_vector(7 downto 0) := "00000011";
  constant CCU_DBG_THREAD_FINISH : std_logic_vector(7 downto 0) := "00000101";
  constant CCU_DBG_WRITE_WP_HIT : std_logic_vector(7 downto 0) := "00000100";
  constant CCU_TEU_CLEAR_BP : std_logic_vector(2 downto 0) := "010";
  constant CCU_TEU_CLEAR_WP : std_logic_vector(2 downto 0) := "100";
  constant CCU_TEU_INTR : std_logic_vector(2 downto 0) := "101";
  constant CCU_TEU_SET_BP : std_logic_vector(2 downto 0) := "001";
  constant CCU_TEU_SET_WP : std_logic_vector(2 downto 0) := "011";
  constant CONTROL_TRANSFER_INSTR : std_logic_vector(2 downto 0) := "011";
  constant CP_DISABLED_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000010000000000000";
  constant CP_DISABLED_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000001100";
  constant CP_EXCEPTION_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000010000000000000000000";
  constant CP_EXCEPTION_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000010010";
  constant CP_INSTR : std_logic_vector(2 downto 0) := "110";
  constant DATA_ACCESS_ERROR_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000100000000000000000000";
  constant DATA_ACCESS_ERROR_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000010011";
  constant DATA_ACCESS_EXCEPTION_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000001000000000000000000000";
  constant DATA_ACCESS_EXCEPTION_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000010100";
  constant DATA_STORE_ERROR_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000000000000100000";
  constant DATA_STORE_ERROR_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000000101";
  constant DATA_TRANSFER_INSTR : std_logic_vector(2 downto 0) := "001";
  constant DEBUG_MODE_MASK : std_logic_vector(7 downto 0) := "00000010";
  constant DIVISION_BY_ZERO_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000100000000000000000000000";
  constant DIVISION_BY_ZERO_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000010110";
  constant EXCEPTION_FOUND : std_logic_vector(7 downto 0) := "00000010";
  constant FOUR_3 : std_logic_vector(2 downto 0) := "100";
  constant FP_DISABLED_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000001000000000000";
  constant FP_DISABLED_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000001011";
  constant FP_EXCEPTION_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000001000000000000000000";
  constant FP_EXCEPTION_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000010001";
  constant FP_INSTR : std_logic_vector(2 downto 0) := "101";
  constant GDB_DBG_CONNECT : std_logic_vector(7 downto 0) := "00001110";
  constant GDB_DBG_CONTINUE : std_logic_vector(7 downto 0) := "00010000";
  constant GDB_DBG_DETACH : std_logic_vector(7 downto 0) := "00001111";
  constant GDB_DBG_KILL : std_logic_vector(7 downto 0) := "00010011";
  constant GDB_DBG_READ_CONTROL_REG : std_logic_vector(7 downto 0) := "00001101";
  constant GDB_DBG_READ_CPUNIT_REG : std_logic_vector(7 downto 0) := "00010001";
  constant GDB_DBG_READ_FPUNIT_REG : std_logic_vector(7 downto 0) := "00000011";
  constant GDB_DBG_READ_INIT_NPC : std_logic_vector(7 downto 0) := "00011101";
  constant GDB_DBG_READ_INIT_PC : std_logic_vector(7 downto 0) := "00011100";
  constant GDB_DBG_READ_INIT_PSR : std_logic_vector(7 downto 0) := "00011110";
  constant GDB_DBG_READ_IUNIT_REG : std_logic_vector(7 downto 0) := "00000001";
  constant GDB_DBG_READ_MEM : std_logic_vector(7 downto 0) := "00000110";
  constant GDB_DBG_READ_MODE : std_logic_vector(7 downto 0) := "00011111";
  constant GDB_DBG_REMOVE_BREAK_POINT : std_logic_vector(7 downto 0) := "00001001";
  constant GDB_DBG_REMOVE_WATCH_POINT : std_logic_vector(7 downto 0) := "00001011";
  constant GDB_DBG_SET_BREAK_POINT : std_logic_vector(7 downto 0) := "00001000";
  constant GDB_DBG_SET_WATCH_POINT : std_logic_vector(7 downto 0) := "00001010";
  constant GDB_DBG_WRITE_CONTROL_REG : std_logic_vector(7 downto 0) := "00010100";
  constant GDB_DBG_WRITE_CPUNIT_REG : std_logic_vector(7 downto 0) := "00010010";
  constant GDB_DBG_WRITE_FPUNIT_REG : std_logic_vector(7 downto 0) := "00000100";
  constant GDB_DBG_WRITE_INIT_NPC : std_logic_vector(7 downto 0) := "00011010";
  constant GDB_DBG_WRITE_INIT_PC : std_logic_vector(7 downto 0) := "00011001";
  constant GDB_DBG_WRITE_INIT_PSR : std_logic_vector(7 downto 0) := "00011011";
  constant GDB_DBG_WRITE_IUNIT_REG : std_logic_vector(7 downto 0) := "00000010";
  constant GDB_DBG_WRITE_MEM : std_logic_vector(7 downto 0) := "00000111";
  constant GDB_DBG_WRITE_RESET : std_logic_vector(7 downto 0) := "00011000";
  constant HARDWARE_ERROR_TRAP_BIT_VEC : std_logic_vector(7 downto 0) := "00100000";
  constant HARDWARE_ERROR_TRAP_INDEX : std_logic_vector(7 downto 0) := "00000101";
  constant HARD_RESET_MASK : std_logic_vector(7 downto 0) := "00000001";
  constant IEEE_754_EXCEPTION_TRAP_BIT_VEC : std_logic_vector(7 downto 0) := "00000010";
  constant IEEE_754_EXCEPTION_TRAP_INDEX : std_logic_vector(7 downto 0) := "00000001";
  constant ILLEGAL_INSTR : std_logic_vector(2 downto 0) := "111";
  constant ILLEGAL_INSTRUCTION_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000000010000000000";
  constant ILLEGAL_INSTRUCTION_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000001001";
  constant ILLEGAL_IU_INSTRUCTION_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000000100000000000";
  constant ILLEGAL_IU_INSTRUCTION_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000001010";
  constant INIT_ASR_AND_WINDOW_REGS : std_logic_vector(2 downto 0) := "111";
  constant INSTRUCTION_ACCESS_ERROR_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000000000010000000";
  constant INSTRUCTION_ACCESS_ERROR_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000000110";
  constant INSTRUCTION_ACCESS_EXCEPTION_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000000000000010000";
  constant INSTRUCTION_ACCESS_EXCEPTION_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000000100";
  constant INTERRUPT_FOUND : std_logic_vector(7 downto 0) := "00000001";
  constant INVALID_FP_REGISTER_TRAP_BIT_VEC : std_logic_vector(7 downto 0) := "01000000";
  constant INVALID_FP_REGISTER_TRAP_INDEX : std_logic_vector(7 downto 0) := "00000110";
  constant KILL_STREAM_MASK : std_logic_vector(7 downto 0) := "10000000";
  constant KILL_THREAD_MASK : std_logic_vector(7 downto 0) := "10000000";
  constant LOGGER_ACTIVE_MASK : std_logic_vector(7 downto 0) := "00001000";
  constant MACHINE_ERROR : std_logic_vector(7 downto 0) := "00000011";
  constant MAE_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000000000000000100";
  constant MAE_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000000010";
  constant MEM_ADDRESS_NOT_ALIGNED_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000100000000000000000";
  constant MEM_ADDRESS_NOT_ALIGNED_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000010000";
  constant MISC_INSTR : std_logic_vector(2 downto 0) := "100";
  constant MMU_PASS_THROUGH_HLIMIT : std_logic_vector(7 downto 0) := "00101111";
  constant MMU_PASS_THROUGH_LLIMIT : std_logic_vector(7 downto 0) := "00100000";
  constant MMU_READ_DWORD : std_logic_vector(7 downto 0) := "00000010";
  constant MMU_READ_LINE : std_logic_vector(7 downto 0) := "00000011";
  constant MMU_WRITE_DWORD : std_logic_vector(7 downto 0) := "00000001";
  constant MMU_WRITE_DWORD_AND_READ_LINE : std_logic_vector(7 downto 0) := "00000111";
  constant MMU_WRITE_DWORD_NO_RESPONSE : std_logic_vector(7 downto 0) := "00000101";
  constant MMU_WRITE_FSR : std_logic_vector(7 downto 0) := "00000100";
  constant NEW_STREAM_MASK : std_logic_vector(7 downto 0) := "10000000";
  constant NEW_THREAD_MASK : std_logic_vector(7 downto 0) := "10000000";
  constant NONE_TRAP_BIT_VEC : std_logic_vector(7 downto 0) := "00000001";
  constant NONE_TRAP_INDEX : std_logic_vector(7 downto 0) := "00000000";
  constant NOP_INSTRUCTION : std_logic_vector(31 downto 0) := "00000001000000000000000000000000";
  constant NO_BLOCK_READ : std_logic_vector(0 downto 0) := "0";
  constant NPC_RESET_VALUE : std_logic_vector(31 downto 0) := "00000000000000000000000000000100";
  constant NWINDOWS : std_logic_vector(31 downto 0) := "00000000000000000000000000001000";
  constant NWINDOWS_MOD_MASK_32 : std_logic_vector(31 downto 0) := "00000000000000000000000000000111";
  constant NWINDOWS_MOD_MASK_5 : std_logic_vector(4 downto 0) := "00111";
  constant NWINDOWSx16 : std_logic_vector(31 downto 0) := "00000000000000000000000010000000";
  constant NWINDOWSx16_MOD_MASK_32 : std_logic_vector(31 downto 0) := "00000000000000000000000001111111";
  constant NWINDOWSx2 : std_logic_vector(31 downto 0) := "00000000000000000000000000010000";
  constant ONE_1 : std_logic_vector(0 downto 0) := "1";
  constant ONE_10 : std_logic_vector(9 downto 0) := "0000000001";
  constant ONE_11 : std_logic_vector(10 downto 0) := "00000000001";
  constant ONE_12 : std_logic_vector(11 downto 0) := "000000000001";
  constant ONE_128 : std_logic_vector(127 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
  constant ONE_13 : std_logic_vector(12 downto 0) := "0000000000001";
  constant ONE_14 : std_logic_vector(13 downto 0) := "00000000000001";
  constant ONE_16 : std_logic_vector(15 downto 0) := "0000000000000001";
  constant ONE_17 : std_logic_vector(16 downto 0) := "00000000000000001";
  constant ONE_18 : std_logic_vector(17 downto 0) := "000000000000000001";
  constant ONE_19 : std_logic_vector(18 downto 0) := "0000000000000000001";
  constant ONE_2 : std_logic_vector(1 downto 0) := "01";
  constant ONE_20 : std_logic_vector(19 downto 0) := "00000000000000000001";
  constant ONE_23 : std_logic_vector(22 downto 0) := "00000000000000000000001";
  constant ONE_24 : std_logic_vector(23 downto 0) := "000000000000000000000001";
  constant ONE_25 : std_logic_vector(24 downto 0) := "0000000000000000000000001";
  constant ONE_256 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
  constant ONE_29 : std_logic_vector(28 downto 0) := "00000000000000000000000000001";
  constant ONE_3 : std_logic_vector(2 downto 0) := "001";
  constant ONE_31 : std_logic_vector(30 downto 0) := "0000000000000000000000000000001";
  constant ONE_32 : std_logic_vector(31 downto 0) := "00000000000000000000000000000001";
  constant ONE_36 : std_logic_vector(35 downto 0) := "000000000000000000000000000000000001";
  constant ONE_4 : std_logic_vector(3 downto 0) := "0001";
  constant ONE_48 : std_logic_vector(47 downto 0) := "000000000000000000000000000000000000000000000001";
  constant ONE_5 : std_logic_vector(4 downto 0) := "00001";
  constant ONE_52 : std_logic_vector(51 downto 0) := "0000000000000000000000000000000000000000000000000001";
  constant ONE_6 : std_logic_vector(5 downto 0) := "000001";
  constant ONE_62 : std_logic_vector(61 downto 0) := "00000000000000000000000000000000000000000000000000000000000001";
  constant ONE_63 : std_logic_vector(62 downto 0) := "000000000000000000000000000000000000000000000000000000000000001";
  constant ONE_64 : std_logic_vector(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000001";
  constant ONE_7 : std_logic_vector(6 downto 0) := "0000001";
  constant ONE_8 : std_logic_vector(7 downto 0) := "00000001";
  constant ONE_9 : std_logic_vector(8 downto 0) := "000000001";
  constant PC_RESET_VALUE : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
  constant PRIVILEGED_INSTRUCTION_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000000001000000000";
  constant PRIVILEGED_INSTRUCTION_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000001000";
  constant PROCESSOR_ERROR_MODE : std_logic_vector(1 downto 0) := "11";
  constant PROCESSOR_EXECUTE_MODE : std_logic_vector(1 downto 0) := "10";
  constant PROCESSOR_RESET_MODE : std_logic_vector(1 downto 0) := "01";
  constant PROCESSOR_UNDEFINED_MODE : std_logic_vector(1 downto 0) := "00";
  constant PSR_RESET_VALUE : std_logic_vector(31 downto 0) := "00000000000000000001000011000000";
  constant REQUEST_TYPE_BRIDGE_CONFIG_READ : std_logic_vector(3 downto 0) := "1001";
  constant REQUEST_TYPE_BRIDGE_CONFIG_WRITE : std_logic_vector(3 downto 0) := "1000";
  constant REQUEST_TYPE_CCU_CACHE_READ : std_logic_vector(3 downto 0) := "0101";
  constant REQUEST_TYPE_CCU_CACHE_WRITE : std_logic_vector(3 downto 0) := "0110";
  constant REQUEST_TYPE_IFETCH : std_logic_vector(3 downto 0) := "0000";
  constant REQUEST_TYPE_NOP : std_logic_vector(3 downto 0) := "0111";
  constant REQUEST_TYPE_READ : std_logic_vector(3 downto 0) := "0001";
  constant REQUEST_TYPE_STBAR : std_logic_vector(3 downto 0) := "0011";
  constant REQUEST_TYPE_WRFSRFAR : std_logic_vector(3 downto 0) := "0100";
  constant REQUEST_TYPE_WRITE : std_logic_vector(3 downto 0) := "0010";
  constant RESERVED_TRAP_BIT_VEC : std_logic_vector(7 downto 0) := "10000000";
  constant RESERVED_TRAP_INDEX : std_logic_vector(7 downto 0) := "00000111";
  constant RESET_TRAP_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000000000000000010";
  constant RESET_TRAP_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000000001";
  constant R_REGISTER_ACCESS_ERROR_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000000000100000000";
  constant R_REGISTER_ACCESS_ERROR_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000000111";
  constant SEQUENCE_ERROR_TRAP_BIT_VEC : std_logic_vector(7 downto 0) := "00010000";
  constant SEQUENCE_ERROR_TRAP_INDEX : std_logic_vector(7 downto 0) := "00000100";
  constant SINGLE_STEP_MASK : std_logic_vector(7 downto 0) := "00000100";
  constant TAG_OVERFLOW_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000010000000000000000000000";
  constant TAG_OVERFLOW_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000010101";
  constant TEU_ANNUL_NEXT_INDEX : std_logic_vector(7 downto 0) := "00000110";
  constant TEU_DBG_BREAK_POINT_INDEX : std_logic_vector(7 downto 0) := "00000011";
  constant TEU_DBG_WATCH_POINT_INDEX : std_logic_vector(7 downto 0) := "00000100";
  constant TEU_EXCEPTION_INDEX : std_logic_vector(7 downto 0) := "00000010";
  constant TEU_FETCH_IS_SPINNING : std_logic_vector(7 downto 0) := "00000111";
  constant TEU_INTERRUPT_INDEX : std_logic_vector(7 downto 0) := "00000001";
  constant TEU_MACHINE_ERROR_INDEX : std_logic_vector(7 downto 0) := "00000000";
  constant TEU_SINGLE_STEP_INDEX : std_logic_vector(7 downto 0) := "00000101";
  constant THREE_2 : std_logic_vector(1 downto 0) := "11";
  constant THREE_3 : std_logic_vector(2 downto 0) := "011";
  constant TRACE_ON : std_logic_vector(0 downto 0) := "1";
  constant TRAP_INSTRUCTION_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000001000000000000000000000000";
  constant TRAP_INSTRUCTION_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000010111";
  constant TRAP_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000000000000000001";
  constant TRAP_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
  constant TT_MASK : std_logic_vector(31 downto 0) := "11111111111111111111000000001111";
  constant TWO_2 : std_logic_vector(1 downto 0) := "10";
  constant TWO_3 : std_logic_vector(2 downto 0) := "010";
  constant UNFINISHED_FPOP_TRAP_BIT_VEC : std_logic_vector(7 downto 0) := "00000100";
  constant UNFINISHED_FPOP_TRAP_INDEX : std_logic_vector(7 downto 0) := "00000010";
  constant UNIMPLEMENTED_FLUSH_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000000100000000000000";
  constant UNIMPLEMENTED_FLUSH_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000001101";
  constant UNIMPLEMENTED_FPOP_TRAP_BIT_VEC : std_logic_vector(7 downto 0) := "00001000";
  constant UNIMPLEMENTED_FPOP_TRAP_INDEX : std_logic_vector(7 downto 0) := "00000011";
  constant WIM_MASK : std_logic_vector(31 downto 0) := "00000000000000000000000011111111";
  constant WINDOW_OVERFLOW_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000001000000000000000";
  constant WINDOW_OVERFLOW_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000001110";
  constant WINDOW_UNDERFLOW_TRAP_BIT_VEC : std_logic_vector(31 downto 0) := "00000000000000010000000000000000";
  constant WINDOW_UNDERFLOW_TRAP_INDEX : std_logic_vector(31 downto 0) := "00000000000000000000000000001111";
  constant ZERO_1 : std_logic_vector(0 downto 0) := "0";
  constant ZERO_10 : std_logic_vector(9 downto 0) := "0000000000";
  constant ZERO_11 : std_logic_vector(10 downto 0) := "00000000000";
  constant ZERO_12 : std_logic_vector(11 downto 0) := "000000000000";
  constant ZERO_128 : std_logic_vector(127 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant ZERO_13 : std_logic_vector(12 downto 0) := "0000000000000";
  constant ZERO_14 : std_logic_vector(13 downto 0) := "00000000000000";
  constant ZERO_16 : std_logic_vector(15 downto 0) := "0000000000000000";
  constant ZERO_17 : std_logic_vector(16 downto 0) := "00000000000000000";
  constant ZERO_18 : std_logic_vector(17 downto 0) := "000000000000000000";
  constant ZERO_19 : std_logic_vector(18 downto 0) := "0000000000000000000";
  constant ZERO_2 : std_logic_vector(1 downto 0) := "00";
  constant ZERO_20 : std_logic_vector(19 downto 0) := "00000000000000000000";
  constant ZERO_23 : std_logic_vector(22 downto 0) := "00000000000000000000000";
  constant ZERO_24 : std_logic_vector(23 downto 0) := "000000000000000000000000";
  constant ZERO_25 : std_logic_vector(24 downto 0) := "0000000000000000000000000";
  constant ZERO_256 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant ZERO_29 : std_logic_vector(28 downto 0) := "00000000000000000000000000000";
  constant ZERO_3 : std_logic_vector(2 downto 0) := "000";
  constant ZERO_31 : std_logic_vector(30 downto 0) := "0000000000000000000000000000000";
  constant ZERO_32 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
  constant ZERO_36 : std_logic_vector(35 downto 0) := "000000000000000000000000000000000000";
  constant ZERO_4 : std_logic_vector(3 downto 0) := "0000";
  constant ZERO_48 : std_logic_vector(47 downto 0) := "000000000000000000000000000000000000000000000000";
  constant ZERO_5 : std_logic_vector(4 downto 0) := "00000";
  constant ZERO_52 : std_logic_vector(51 downto 0) := "0000000000000000000000000000000000000000000000000000";
  constant ZERO_6 : std_logic_vector(5 downto 0) := "000000";
  constant ZERO_62 : std_logic_vector(61 downto 0) := "00000000000000000000000000000000000000000000000000000000000000";
  constant ZERO_63 : std_logic_vector(62 downto 0) := "000000000000000000000000000000000000000000000000000000000000000";
  constant ZERO_64 : std_logic_vector(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000";
  constant ZERO_7 : std_logic_vector(6 downto 0) := "0000000";
  constant ZERO_8 : std_logic_vector(7 downto 0) := "00000000";
  constant ZERO_9 : std_logic_vector(8 downto 0) := "000000000";
  constant default_mem_pool_base_address : std_logic_vector(0 downto 0) := "0";
  component iu_exec is -- 
    port (-- 
      clk : in std_logic;
      reset : in std_logic;
      iunit_exec_fast_alu_result_to_writeback_pipe_read_data: out std_logic_vector(108 downto 0);
      iunit_exec_fast_alu_result_to_writeback_pipe_read_req : in std_logic_vector(0 downto 0);
      iunit_exec_fast_alu_result_to_writeback_pipe_read_ack : out std_logic_vector(0 downto 0);
      iunit_exec_to_writeback_pipe_read_data: out std_logic_vector(125 downto 0);
      iunit_exec_to_writeback_pipe_read_req : in std_logic_vector(0 downto 0);
      iunit_exec_to_writeback_pipe_read_ack : out std_logic_vector(0 downto 0);
      iunit_register_file_read_access_response_pipe_write_data: in std_logic_vector(141 downto 0);
      iunit_register_file_read_access_response_pipe_write_req : in std_logic_vector(0 downto 0);
      iunit_register_file_read_access_response_pipe_write_ack : out std_logic_vector(0 downto 0);
      noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_read_data: out std_logic_vector(16 downto 0);
      noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_read_req : in std_logic_vector(0 downto 0);
      noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_read_ack : out std_logic_vector(0 downto 0);
      noblock_iunit_exec_bypass_signal_to_register_file_pipe_read_data: out std_logic_vector(82 downto 0);
      noblock_iunit_exec_bypass_signal_to_register_file_pipe_read_req : in std_logic_vector(0 downto 0);
      noblock_iunit_exec_bypass_signal_to_register_file_pipe_read_ack : out std_logic_vector(0 downto 0);
      noblock_iunit_exec_to_regfile_credit_return_pipe_read_data: out std_logic_vector(0 downto 0);
      noblock_iunit_exec_to_regfile_credit_return_pipe_read_req : in std_logic_vector(0 downto 0);
      noblock_iunit_exec_to_regfile_credit_return_pipe_read_ack : out std_logic_vector(0 downto 0);
      teu_idispatch_to_iunit_exec_pipe_write_data: in std_logic_vector(149 downto 0);
      teu_idispatch_to_iunit_exec_pipe_write_req : in std_logic_vector(0 downto 0);
      teu_idispatch_to_iunit_exec_pipe_write_ack : out std_logic_vector(0 downto 0);
      teu_iunit_to_stream_corrector_pipe_read_data: out std_logic_vector(89 downto 0);
      teu_iunit_to_stream_corrector_pipe_read_req : in std_logic_vector(0 downto 0);
      teu_iunit_to_stream_corrector_pipe_read_ack : out std_logic_vector(0 downto 0);
      teu_iunit_trap_to_fpunit_pipe_read_data: out std_logic_vector(12 downto 0);
      teu_iunit_trap_to_fpunit_pipe_read_req : in std_logic_vector(0 downto 0);
      teu_iunit_trap_to_fpunit_pipe_read_ack : out std_logic_vector(0 downto 0);
      teu_iunit_trap_to_loadstore_pipe_read_data: out std_logic_vector(0 downto 0);
      teu_iunit_trap_to_loadstore_pipe_read_req : in std_logic_vector(0 downto 0);
      teu_iunit_trap_to_loadstore_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
    -- 
  end component;
  -- 
end package iu_exec_global_package;
-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity alignDivisorToDividendRevised_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    DIVIDEND : in  std_logic_vector(63 downto 0);
    udivisor : in  std_logic_vector(31 downto 0);
    SHIFTED_DIVIDEND : out  std_logic_vector(63 downto 0);
    SHIFTED_DIVISOR : out  std_logic_vector(31 downto 0);
    INITIAL_QMASK : out  std_logic_vector(63 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity alignDivisorToDividendRevised_Operator;
architecture alignDivisorToDividendRevised_Operator_arch of alignDivisorToDividendRevised_Operator is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal update_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal DIVIDEND_buffer :  std_logic_vector(63 downto 0);
  signal DIVIDEND_update_enable: Boolean;
  signal DIVIDEND_update_enable_unmarked: Boolean;
  signal udivisor_buffer :  std_logic_vector(31 downto 0);
  signal udivisor_update_enable: Boolean;
  signal udivisor_update_enable_unmarked: Boolean;
  -- output port buffer signals
  signal SHIFTED_DIVIDEND_buffer :  std_logic_vector(63 downto 0);
  signal SHIFTED_DIVIDEND_update_enable: Boolean;
  signal SHIFTED_DIVISOR_buffer :  std_logic_vector(31 downto 0);
  signal SHIFTED_DIVISOR_update_enable: Boolean;
  signal INITIAL_QMASK_buffer :  std_logic_vector(63 downto 0);
  signal INITIAL_QMASK_update_enable: Boolean;
  signal alignDivisorToDividendRevised_CP_138_start: Boolean;
  signal alignDivisorToDividendRevised_CP_138_symbol: Boolean;
  signal cp_all_inputs_sampled: Boolean;
  -- volatile/operator module components. 
  component u_set_index_64_Volatile is -- 
    port ( -- 
      idx : in  std_logic_vector(5 downto 0);
      x : out  std_logic_vector(63 downto 0)-- 
    );
    -- 
  end component; 
  component find_left_32_Volatile is -- 
    port ( -- 
      fp_32 : in  std_logic_vector(31 downto 0);
      position : out  std_logic_vector(4 downto 0);
      found : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component find_leftmost_64_Volatile is -- 
    port ( -- 
      fp_64 : in  std_logic_vector(63 downto 0);
      position : out  std_logic_vector(5 downto 0);
      found : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component u64_sll_Volatile is -- 
    port ( -- 
      X : in  std_logic_vector(63 downto 0);
      S : in  std_logic_vector(6 downto 0);
      Y : out  std_logic_vector(63 downto 0)-- 
    );
    -- 
  end component; 
  component u32_sll_Volatile is -- 
    port ( -- 
      X : in  std_logic_vector(31 downto 0);
      S : in  std_logic_vector(5 downto 0);
      Y : out  std_logic_vector(31 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal W_INITIAL_QMASK_1655_inst_req_0 : boolean;
  signal W_INITIAL_QMASK_1655_inst_ack_0 : boolean;
  signal W_INITIAL_QMASK_1655_inst_req_1 : boolean;
  signal W_INITIAL_QMASK_1655_inst_ack_1 : boolean;
  signal W_SHIFTED_DIVISOR_1658_inst_req_0 : boolean;
  signal W_SHIFTED_DIVISOR_1658_inst_ack_0 : boolean;
  signal W_SHIFTED_DIVISOR_1658_inst_req_1 : boolean;
  signal W_SHIFTED_DIVISOR_1658_inst_ack_1 : boolean;
  signal W_SHIFTED_DIVIDEND_1661_inst_req_0 : boolean;
  signal W_SHIFTED_DIVIDEND_1661_inst_ack_0 : boolean;
  signal W_SHIFTED_DIVIDEND_1661_inst_req_1 : boolean;
  signal W_SHIFTED_DIVIDEND_1661_inst_ack_1 : boolean;
  -- 
begin --  
  -- sample-ack is join of  cp-entry-symbol and all-inputs-sampled 
  sample_ack <= cp_all_inputs_sampled;
  -- input handling ------------------------------------------------
  DIVIDEND_buffer <= DIVIDEND;
  udivisor_buffer <= udivisor;
  -- join of sample-req and update-ack-symbol.. used to trigger CP.
  alignDivisorToDividendRevised_CP_138_start_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 3);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 3);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 47) := "alignDivisorToDividendRevised_CP_138_start_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sample_req & update_ack_symbol;
    gj_alignDivisorToDividendRevised_CP_138_start_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => alignDivisorToDividendRevised_CP_138_start, clk => clk, reset => reset); --
  end block;
  -- join of all input-sampled signals.. used to produce sample_ack.
  cp_all_inputs_sampled_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
    constant joinName: string(1 to 26) := "cp_all_inputs_sampled_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= DIVIDEND_update_enable_unmarked & udivisor_update_enable_unmarked;
    gj_cp_all_inputs_sampled_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => cp_all_inputs_sampled, clk => clk, reset => reset); --
  end block;
  -- output handling  -------------------------------------------------------
  SHIFTED_DIVIDEND <= SHIFTED_DIVIDEND_buffer;
  SHIFTED_DIVIDEND_update_enable <= update_req;
  SHIFTED_DIVISOR <= SHIFTED_DIVISOR_buffer;
  SHIFTED_DIVISOR_update_enable <= update_req;
  INITIAL_QMASK <= INITIAL_QMASK_buffer;
  INITIAL_QMASK_update_enable <= update_req;
  update_ack_symbol <= alignDivisorToDividendRevised_CP_138_symbol;
  update_ack <= update_ack_symbol;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  alignDivisorToDividendRevised_CP_138: Block -- control-path 
    signal alignDivisorToDividendRevised_CP_138_elements: BooleanArray(29 downto 0);
    -- 
  begin -- 
    alignDivisorToDividendRevised_CP_138_elements(0) <= alignDivisorToDividendRevised_CP_138_start;
    alignDivisorToDividendRevised_CP_138_symbol <= alignDivisorToDividendRevised_CP_138_elements(29);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	13 
    -- CP-element group 1: 	9 
    -- CP-element group 1: 	17 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_1620_to_assign_stmt_1663/$entry
      -- 
    alignDivisorToDividendRevised_CP_138_elements(1) <= alignDivisorToDividendRevised_CP_138_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	19 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	22 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_1620_to_assign_stmt_1663/DIVIDEND_update_enable
      -- CP-element group 2: 	 call_stmt_1620_to_assign_stmt_1663/DIVIDEND_update_enable_out
      -- 
    alignDivisorToDividendRevised_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 48) := "alignDivisorToDividendRevised_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= alignDivisorToDividendRevised_CP_138_elements(11) & alignDivisorToDividendRevised_CP_138_elements(19);
      gj_alignDivisorToDividendRevised_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => alignDivisorToDividendRevised_CP_138_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	11 
    -- CP-element group 3: 	19 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	23 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_1620_to_assign_stmt_1663/DIVIDEND_update_enable_unmarked
      -- CP-element group 3: 	 call_stmt_1620_to_assign_stmt_1663/DIVIDEND_update_enable_unmarked_out
      -- 
    alignDivisorToDividendRevised_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 48) := "alignDivisorToDividendRevised_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= alignDivisorToDividendRevised_CP_138_elements(11) & alignDivisorToDividendRevised_CP_138_elements(19);
      gj_alignDivisorToDividendRevised_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => alignDivisorToDividendRevised_CP_138_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	11 
    -- CP-element group 4: 	15 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	24 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 call_stmt_1620_to_assign_stmt_1663/udivisor_update_enable
      -- CP-element group 4: 	 call_stmt_1620_to_assign_stmt_1663/udivisor_update_enable_out
      -- 
    alignDivisorToDividendRevised_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 48) := "alignDivisorToDividendRevised_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= alignDivisorToDividendRevised_CP_138_elements(11) & alignDivisorToDividendRevised_CP_138_elements(15);
      gj_alignDivisorToDividendRevised_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => alignDivisorToDividendRevised_CP_138_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	11 
    -- CP-element group 5: 	15 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	25 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 call_stmt_1620_to_assign_stmt_1663/udivisor_update_enable_unmarked
      -- CP-element group 5: 	 call_stmt_1620_to_assign_stmt_1663/udivisor_update_enable_unmarked_out
      -- 
    alignDivisorToDividendRevised_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 48) := "alignDivisorToDividendRevised_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= alignDivisorToDividendRevised_CP_138_elements(11) & alignDivisorToDividendRevised_CP_138_elements(15);
      gj_alignDivisorToDividendRevised_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => alignDivisorToDividendRevised_CP_138_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	26 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	18 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 call_stmt_1620_to_assign_stmt_1663/SHIFTED_DIVIDEND_update_enable
      -- CP-element group 6: 	 call_stmt_1620_to_assign_stmt_1663/SHIFTED_DIVIDEND_update_enable_in
      -- 
    alignDivisorToDividendRevised_CP_138_elements(6) <= alignDivisorToDividendRevised_CP_138_elements(26);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	27 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	14 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 call_stmt_1620_to_assign_stmt_1663/SHIFTED_DIVISOR_update_enable
      -- CP-element group 7: 	 call_stmt_1620_to_assign_stmt_1663/SHIFTED_DIVISOR_update_enable_in
      -- 
    alignDivisorToDividendRevised_CP_138_elements(7) <= alignDivisorToDividendRevised_CP_138_elements(27);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	28 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 call_stmt_1620_to_assign_stmt_1663/INITIAL_QMASK_update_enable
      -- CP-element group 8: 	 call_stmt_1620_to_assign_stmt_1663/INITIAL_QMASK_update_enable_in
      -- 
    alignDivisorToDividendRevised_CP_138_elements(8) <= alignDivisorToDividendRevised_CP_138_elements(28);
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1657_sample_start_
      -- CP-element group 9: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1657_Sample/$entry
      -- CP-element group 9: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1657_Sample/req
      -- 
    req_165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => alignDivisorToDividendRevised_CP_138_elements(9), ack => W_INITIAL_QMASK_1655_inst_req_0); -- 
    alignDivisorToDividendRevised_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 48) := "alignDivisorToDividendRevised_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= alignDivisorToDividendRevised_CP_138_elements(1) & alignDivisorToDividendRevised_CP_138_elements(11);
      gj_alignDivisorToDividendRevised_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => alignDivisorToDividendRevised_CP_138_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1657_update_start_
      -- CP-element group 10: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1657_Update/$entry
      -- CP-element group 10: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1657_Update/req
      -- 
    req_170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => alignDivisorToDividendRevised_CP_138_elements(10), ack => W_INITIAL_QMASK_1655_inst_req_1); -- 
    alignDivisorToDividendRevised_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "alignDivisorToDividendRevised_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= alignDivisorToDividendRevised_CP_138_elements(8) & alignDivisorToDividendRevised_CP_138_elements(12);
      gj_alignDivisorToDividendRevised_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => alignDivisorToDividendRevised_CP_138_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	3 
    -- CP-element group 11: 	5 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	4 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	2 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1657_sample_completed_
      -- CP-element group 11: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1657_Sample/$exit
      -- CP-element group 11: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1657_Sample/ack
      -- 
    ack_166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_INITIAL_QMASK_1655_inst_ack_0, ack => alignDivisorToDividendRevised_CP_138_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	21 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1657_update_completed_
      -- CP-element group 12: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1657_Update/$exit
      -- CP-element group 12: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1657_Update/ack
      -- 
    ack_171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_INITIAL_QMASK_1655_inst_ack_1, ack => alignDivisorToDividendRevised_CP_138_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	1 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1660_sample_start_
      -- CP-element group 13: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1660_Sample/$entry
      -- CP-element group 13: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1660_Sample/req
      -- 
    req_179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => alignDivisorToDividendRevised_CP_138_elements(13), ack => W_SHIFTED_DIVISOR_1658_inst_req_0); -- 
    alignDivisorToDividendRevised_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "alignDivisorToDividendRevised_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= alignDivisorToDividendRevised_CP_138_elements(1) & alignDivisorToDividendRevised_CP_138_elements(15);
      gj_alignDivisorToDividendRevised_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => alignDivisorToDividendRevised_CP_138_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	7 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1660_update_start_
      -- CP-element group 14: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1660_Update/$entry
      -- CP-element group 14: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1660_Update/req
      -- 
    req_184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => alignDivisorToDividendRevised_CP_138_elements(14), ack => W_SHIFTED_DIVISOR_1658_inst_req_1); -- 
    alignDivisorToDividendRevised_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "alignDivisorToDividendRevised_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= alignDivisorToDividendRevised_CP_138_elements(7) & alignDivisorToDividendRevised_CP_138_elements(16);
      gj_alignDivisorToDividendRevised_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => alignDivisorToDividendRevised_CP_138_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	5 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	4 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1660_sample_completed_
      -- CP-element group 15: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1660_Sample/$exit
      -- CP-element group 15: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1660_Sample/ack
      -- 
    ack_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_SHIFTED_DIVISOR_1658_inst_ack_0, ack => alignDivisorToDividendRevised_CP_138_elements(15)); -- 
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1660_update_completed_
      -- CP-element group 16: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1660_Update/$exit
      -- CP-element group 16: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1660_Update/ack
      -- 
    ack_185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_SHIFTED_DIVISOR_1658_inst_ack_1, ack => alignDivisorToDividendRevised_CP_138_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	1 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1663_sample_start_
      -- CP-element group 17: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1663_Sample/$entry
      -- CP-element group 17: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1663_Sample/req
      -- 
    req_193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => alignDivisorToDividendRevised_CP_138_elements(17), ack => W_SHIFTED_DIVIDEND_1661_inst_req_0); -- 
    alignDivisorToDividendRevised_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "alignDivisorToDividendRevised_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= alignDivisorToDividendRevised_CP_138_elements(1) & alignDivisorToDividendRevised_CP_138_elements(19);
      gj_alignDivisorToDividendRevised_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => alignDivisorToDividendRevised_CP_138_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	6 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1663_update_start_
      -- CP-element group 18: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1663_Update/$entry
      -- CP-element group 18: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1663_Update/req
      -- 
    req_198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => alignDivisorToDividendRevised_CP_138_elements(18), ack => W_SHIFTED_DIVIDEND_1661_inst_req_1); -- 
    alignDivisorToDividendRevised_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "alignDivisorToDividendRevised_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= alignDivisorToDividendRevised_CP_138_elements(6) & alignDivisorToDividendRevised_CP_138_elements(20);
      gj_alignDivisorToDividendRevised_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => alignDivisorToDividendRevised_CP_138_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	3 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1663_sample_completed_
      -- CP-element group 19: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1663_Sample/$exit
      -- CP-element group 19: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1663_Sample/ack
      -- 
    ack_194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_SHIFTED_DIVIDEND_1661_inst_ack_0, ack => alignDivisorToDividendRevised_CP_138_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1663_update_completed_
      -- CP-element group 20: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1663_Update/$exit
      -- CP-element group 20: 	 call_stmt_1620_to_assign_stmt_1663/assign_stmt_1663_Update/ack
      -- 
    ack_199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_SHIFTED_DIVIDEND_1661_inst_ack_1, ack => alignDivisorToDividendRevised_CP_138_elements(20)); -- 
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: 	16 
    -- CP-element group 21: 	12 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	29 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 call_stmt_1620_to_assign_stmt_1663/$exit
      -- 
    alignDivisorToDividendRevised_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "alignDivisorToDividendRevised_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= alignDivisorToDividendRevised_CP_138_elements(20) & alignDivisorToDividendRevised_CP_138_elements(16) & alignDivisorToDividendRevised_CP_138_elements(12);
      gj_alignDivisorToDividendRevised_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => alignDivisorToDividendRevised_CP_138_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  place  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 DIVIDEND_update_enable
      -- 
    alignDivisorToDividendRevised_CP_138_elements(22) <= alignDivisorToDividendRevised_CP_138_elements(2);
    -- CP-element group 23:  place  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	3 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 DIVIDEND_update_enable_unmarked
      -- 
    alignDivisorToDividendRevised_CP_138_elements(23) <= alignDivisorToDividendRevised_CP_138_elements(3);
    -- CP-element group 24:  place  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	4 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 udivisor_update_enable
      -- 
    alignDivisorToDividendRevised_CP_138_elements(24) <= alignDivisorToDividendRevised_CP_138_elements(4);
    -- CP-element group 25:  place  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	5 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 udivisor_update_enable_unmarked
      -- 
    alignDivisorToDividendRevised_CP_138_elements(25) <= alignDivisorToDividendRevised_CP_138_elements(5);
    -- CP-element group 26:  place  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	6 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 SHIFTED_DIVIDEND_update_enable
      -- 
    -- CP-element group 27:  place  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	7 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 SHIFTED_DIVISOR_update_enable
      -- 
    -- CP-element group 28:  place  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	8 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 INITIAL_QMASK_update_enable
      -- 
    -- CP-element group 29:  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	21 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 $exit
      -- 
    alignDivisorToDividendRevised_CP_138_elements(29) <= alignDivisorToDividendRevised_CP_138_elements(21);
    --  hookup: inputs to control-path 
    alignDivisorToDividendRevised_CP_138_elements(26) <= SHIFTED_DIVIDEND_update_enable;
    alignDivisorToDividendRevised_CP_138_elements(27) <= SHIFTED_DIVISOR_update_enable;
    alignDivisorToDividendRevised_CP_138_elements(28) <= INITIAL_QMASK_update_enable;
    -- hookup: output from control-path 
    DIVIDEND_update_enable <= alignDivisorToDividendRevised_CP_138_elements(22);
    DIVIDEND_update_enable_unmarked <= alignDivisorToDividendRevised_CP_138_elements(23);
    udivisor_update_enable <= alignDivisorToDividendRevised_CP_138_elements(24);
    udivisor_update_enable_unmarked <= alignDivisorToDividendRevised_CP_138_elements(25);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal SUB_u6_u6_1646_wire : std_logic_vector(5 downto 0);
    signal SUB_u7_u7_1639_wire : std_logic_vector(6 downto 0);
    signal ccq_shift_amount_1651 : std_logic_vector(5 downto 0);
    signal ccq_v_1654 : std_logic_vector(63 downto 0);
    signal konst_1636_wire_constant : std_logic_vector(6 downto 0);
    signal konst_1643_wire_constant : std_logic_vector(5 downto 0);
    signal l_DIVIDEND_1620 : std_logic_vector(5 downto 0);
    signal l_udivisor_1624 : std_logic_vector(4 downto 0);
    signal sdividend_1641 : std_logic_vector(63 downto 0);
    signal sdivisor_1648 : std_logic_vector(31 downto 0);
    signal shift_amount_1634 : std_logic_vector(5 downto 0);
    signal type_cast_1632_wire : std_logic_vector(5 downto 0);
    signal type_cast_1638_wire : std_logic_vector(6 downto 0);
    signal type_cast_1645_wire : std_logic_vector(5 downto 0);
    signal z_DIVIDEND_1620 : std_logic_vector(0 downto 0);
    signal z_udivisor_1624 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_1636_wire_constant <= "0111111";
    konst_1643_wire_constant <= "011111";
    W_INITIAL_QMASK_1655_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_INITIAL_QMASK_1655_inst_req_0;
      W_INITIAL_QMASK_1655_inst_ack_0<= wack(0);
      rreq(0) <= W_INITIAL_QMASK_1655_inst_req_1;
      W_INITIAL_QMASK_1655_inst_ack_1<= rack(0);
      W_INITIAL_QMASK_1655_inst : InterlockBuffer generic map ( -- 
        name => "W_INITIAL_QMASK_1655_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ccq_v_1654,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => INITIAL_QMASK_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_SHIFTED_DIVIDEND_1661_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_SHIFTED_DIVIDEND_1661_inst_req_0;
      W_SHIFTED_DIVIDEND_1661_inst_ack_0<= wack(0);
      rreq(0) <= W_SHIFTED_DIVIDEND_1661_inst_req_1;
      W_SHIFTED_DIVIDEND_1661_inst_ack_1<= rack(0);
      W_SHIFTED_DIVIDEND_1661_inst : InterlockBuffer generic map ( -- 
        name => "W_SHIFTED_DIVIDEND_1661_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sdividend_1641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => SHIFTED_DIVIDEND_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_SHIFTED_DIVISOR_1658_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_SHIFTED_DIVISOR_1658_inst_req_0;
      W_SHIFTED_DIVISOR_1658_inst_ack_0<= wack(0);
      rreq(0) <= W_SHIFTED_DIVISOR_1658_inst_req_1;
      W_SHIFTED_DIVISOR_1658_inst_ack_1<= rack(0);
      W_SHIFTED_DIVISOR_1658_inst : InterlockBuffer generic map ( -- 
        name => "W_SHIFTED_DIVISOR_1658_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sdivisor_1648,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => SHIFTED_DIVISOR_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ccq_shift_amount_1649_inst
    process(shift_amount_1634) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := shift_amount_1634(5 downto 0);
      ccq_shift_amount_1651 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1632_inst
    process(l_udivisor_1624) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 4 downto 0) := l_udivisor_1624(4 downto 0);
      type_cast_1632_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1638_inst
    process(l_DIVIDEND_1620) -- 
      variable tmp_var : std_logic_vector(6 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := l_DIVIDEND_1620(5 downto 0);
      type_cast_1638_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1645_inst
    process(l_udivisor_1624) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 4 downto 0) := l_udivisor_1624(4 downto 0);
      type_cast_1645_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator SUB_u6_u6_1633_inst
    shift_amount_1634 <= std_logic_vector(unsigned(l_DIVIDEND_1620) - unsigned(type_cast_1632_wire));
    -- flow through binary operator SUB_u6_u6_1646_inst
    SUB_u6_u6_1646_wire <= std_logic_vector(unsigned(konst_1643_wire_constant) - unsigned(type_cast_1645_wire));
    -- flow through binary operator SUB_u7_u7_1639_inst
    SUB_u7_u7_1639_wire <= std_logic_vector(unsigned(konst_1636_wire_constant) - unsigned(type_cast_1638_wire));
    volatile_operator_find_leftmost_64_1388: find_leftmost_64_Volatile port map(fp_64 => DIVIDEND_buffer, position => l_DIVIDEND_1620, found => z_DIVIDEND_1620); 
    volatile_operator_find_left_32_1389: find_left_32_Volatile port map(fp_32 => udivisor_buffer, position => l_udivisor_1624, found => z_udivisor_1624); 
    volatile_operator_u64_sll_1394: u64_sll_Volatile port map(X => DIVIDEND_buffer, S => SUB_u7_u7_1639_wire, Y => sdividend_1641); 
    volatile_operator_u32_sll_1397: u32_sll_Volatile port map(X => udivisor_buffer, S => SUB_u6_u6_1646_wire, Y => sdivisor_1648); 
    volatile_operator_u_set_index_64_1399: u_set_index_64_Volatile port map(idx => ccq_shift_amount_1651, x => ccq_v_1654); 
    -- 
  end Block; -- data_path
  -- 
end alignDivisorToDividendRevised_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity decode_alu_exec_control_word_Volatile is -- 
  port ( -- 
    cw : in  std_logic_vector(54 downto 0);
    cti : out  std_logic_vector(0 downto 0);
    is_call : out  std_logic_vector(0 downto 0);
    is_jmpl : out  std_logic_vector(0 downto 0);
    is_rett : out  std_logic_vector(0 downto 0);
    is_bicc : out  std_logic_vector(0 downto 0);
    is_fbfcc : out  std_logic_vector(0 downto 0);
    is_cbccc : out  std_logic_vector(0 downto 0);
    is_ticc : out  std_logic_vector(0 downto 0);
    annul_flag : out  std_logic_vector(0 downto 0);
    br_cond : out  std_logic_vector(3 downto 0);
    alu : out  std_logic_vector(0 downto 0);
    use_alu_add : out  std_logic_vector(0 downto 0);
    is_alu_sub : out  std_logic_vector(0 downto 0);
    is_alu_mul : out  std_logic_vector(0 downto 0);
    is_alu_mulscc : out  std_logic_vector(0 downto 0);
    is_alu_div : out  std_logic_vector(0 downto 0);
    is_alu_sll : out  std_logic_vector(0 downto 0);
    is_alu_srl : out  std_logic_vector(0 downto 0);
    is_alu_sra : out  std_logic_vector(0 downto 0);
    is_alu_and : out  std_logic_vector(0 downto 0);
    is_alu_or : out  std_logic_vector(0 downto 0);
    use_alu_xor : out  std_logic_vector(0 downto 0);
    is_alu_xnor : out  std_logic_vector(0 downto 0);
    signed_mul_div : out  std_logic_vector(0 downto 0);
    negate_second_operand : out  std_logic_vector(0 downto 0);
    with_carry : out  std_logic_vector(0 downto 0);
    set_cc : out  std_logic_vector(0 downto 0);
    tagged_alu_op : out  std_logic_vector(0 downto 0);
    trap_on_overflow : out  std_logic_vector(0 downto 0);
    misc : out  std_logic_vector(0 downto 0);
    is_sethi : out  std_logic_vector(0 downto 0);
    write_psr : out  std_logic_vector(0 downto 0);
    write_wim : out  std_logic_vector(0 downto 0);
    write_tbr : out  std_logic_vector(0 downto 0);
    write_y : out  std_logic_vector(0 downto 0);
    write_asr : out  std_logic_vector(0 downto 0);
    read_psr : out  std_logic_vector(0 downto 0);
    read_wim : out  std_logic_vector(0 downto 0);
    read_tbr : out  std_logic_vector(0 downto 0);
    read_y : out  std_logic_vector(0 downto 0);
    read_asr : out  std_logic_vector(0 downto 0);
    asr_id : out  std_logic_vector(4 downto 0);
    is_save : out  std_logic_vector(0 downto 0);
    is_restore : out  std_logic_vector(0 downto 0);
    dti : out  std_logic_vector(0 downto 0);
    is_iu_dti : out  std_logic_vector(0 downto 0);
    is_load_to_debug : out  std_logic_vector(0 downto 0);
    is_store_to_debug : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity decode_alu_exec_control_word_Volatile;
architecture decode_alu_exec_control_word_Volatile_arch of decode_alu_exec_control_word_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(55-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal cw_buffer :  std_logic_vector(54 downto 0);
  -- output port buffer signals
  signal cti_buffer :  std_logic_vector(0 downto 0);
  signal is_call_buffer :  std_logic_vector(0 downto 0);
  signal is_jmpl_buffer :  std_logic_vector(0 downto 0);
  signal is_rett_buffer :  std_logic_vector(0 downto 0);
  signal is_bicc_buffer :  std_logic_vector(0 downto 0);
  signal is_fbfcc_buffer :  std_logic_vector(0 downto 0);
  signal is_cbccc_buffer :  std_logic_vector(0 downto 0);
  signal is_ticc_buffer :  std_logic_vector(0 downto 0);
  signal annul_flag_buffer :  std_logic_vector(0 downto 0);
  signal br_cond_buffer :  std_logic_vector(3 downto 0);
  signal alu_buffer :  std_logic_vector(0 downto 0);
  signal use_alu_add_buffer :  std_logic_vector(0 downto 0);
  signal is_alu_sub_buffer :  std_logic_vector(0 downto 0);
  signal is_alu_mul_buffer :  std_logic_vector(0 downto 0);
  signal is_alu_mulscc_buffer :  std_logic_vector(0 downto 0);
  signal is_alu_div_buffer :  std_logic_vector(0 downto 0);
  signal is_alu_sll_buffer :  std_logic_vector(0 downto 0);
  signal is_alu_srl_buffer :  std_logic_vector(0 downto 0);
  signal is_alu_sra_buffer :  std_logic_vector(0 downto 0);
  signal is_alu_and_buffer :  std_logic_vector(0 downto 0);
  signal is_alu_or_buffer :  std_logic_vector(0 downto 0);
  signal use_alu_xor_buffer :  std_logic_vector(0 downto 0);
  signal is_alu_xnor_buffer :  std_logic_vector(0 downto 0);
  signal signed_mul_div_buffer :  std_logic_vector(0 downto 0);
  signal negate_second_operand_buffer :  std_logic_vector(0 downto 0);
  signal with_carry_buffer :  std_logic_vector(0 downto 0);
  signal set_cc_buffer :  std_logic_vector(0 downto 0);
  signal tagged_alu_op_buffer :  std_logic_vector(0 downto 0);
  signal trap_on_overflow_buffer :  std_logic_vector(0 downto 0);
  signal misc_buffer :  std_logic_vector(0 downto 0);
  signal is_sethi_buffer :  std_logic_vector(0 downto 0);
  signal write_psr_buffer :  std_logic_vector(0 downto 0);
  signal write_wim_buffer :  std_logic_vector(0 downto 0);
  signal write_tbr_buffer :  std_logic_vector(0 downto 0);
  signal write_y_buffer :  std_logic_vector(0 downto 0);
  signal write_asr_buffer :  std_logic_vector(0 downto 0);
  signal read_psr_buffer :  std_logic_vector(0 downto 0);
  signal read_wim_buffer :  std_logic_vector(0 downto 0);
  signal read_tbr_buffer :  std_logic_vector(0 downto 0);
  signal read_y_buffer :  std_logic_vector(0 downto 0);
  signal read_asr_buffer :  std_logic_vector(0 downto 0);
  signal asr_id_buffer :  std_logic_vector(4 downto 0);
  signal is_save_buffer :  std_logic_vector(0 downto 0);
  signal is_restore_buffer :  std_logic_vector(0 downto 0);
  signal dti_buffer :  std_logic_vector(0 downto 0);
  signal is_iu_dti_buffer :  std_logic_vector(0 downto 0);
  signal is_load_to_debug_buffer :  std_logic_vector(0 downto 0);
  signal is_store_to_debug_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  cw_buffer <= cw;
  -- output handling  -------------------------------------------------------
  cti <= cti_buffer;
  is_call <= is_call_buffer;
  is_jmpl <= is_jmpl_buffer;
  is_rett <= is_rett_buffer;
  is_bicc <= is_bicc_buffer;
  is_fbfcc <= is_fbfcc_buffer;
  is_cbccc <= is_cbccc_buffer;
  is_ticc <= is_ticc_buffer;
  annul_flag <= annul_flag_buffer;
  br_cond <= br_cond_buffer;
  alu <= alu_buffer;
  use_alu_add <= use_alu_add_buffer;
  is_alu_sub <= is_alu_sub_buffer;
  is_alu_mul <= is_alu_mul_buffer;
  is_alu_mulscc <= is_alu_mulscc_buffer;
  is_alu_div <= is_alu_div_buffer;
  is_alu_sll <= is_alu_sll_buffer;
  is_alu_srl <= is_alu_srl_buffer;
  is_alu_sra <= is_alu_sra_buffer;
  is_alu_and <= is_alu_and_buffer;
  is_alu_or <= is_alu_or_buffer;
  use_alu_xor <= use_alu_xor_buffer;
  is_alu_xnor <= is_alu_xnor_buffer;
  signed_mul_div <= signed_mul_div_buffer;
  negate_second_operand <= negate_second_operand_buffer;
  with_carry <= with_carry_buffer;
  set_cc <= set_cc_buffer;
  tagged_alu_op <= tagged_alu_op_buffer;
  trap_on_overflow <= trap_on_overflow_buffer;
  misc <= misc_buffer;
  is_sethi <= is_sethi_buffer;
  write_psr <= write_psr_buffer;
  write_wim <= write_wim_buffer;
  write_tbr <= write_tbr_buffer;
  write_y <= write_y_buffer;
  write_asr <= write_asr_buffer;
  read_psr <= read_psr_buffer;
  read_wim <= read_wim_buffer;
  read_tbr <= read_tbr_buffer;
  read_y <= read_y_buffer;
  read_asr <= read_asr_buffer;
  asr_id <= asr_id_buffer;
  is_save <= is_save_buffer;
  is_restore <= is_restore_buffer;
  dti <= dti_buffer;
  is_iu_dti <= is_iu_dti_buffer;
  is_load_to_debug <= is_load_to_debug_buffer;
  is_store_to_debug <= is_store_to_debug_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- flow-through slice operator slice_2101_inst
    cti_buffer <= cw_buffer(54 downto 54);
    -- flow-through slice operator slice_2105_inst
    is_call_buffer <= cw_buffer(53 downto 53);
    -- flow-through slice operator slice_2109_inst
    is_jmpl_buffer <= cw_buffer(52 downto 52);
    -- flow-through slice operator slice_2113_inst
    is_rett_buffer <= cw_buffer(51 downto 51);
    -- flow-through slice operator slice_2117_inst
    is_bicc_buffer <= cw_buffer(50 downto 50);
    -- flow-through slice operator slice_2121_inst
    is_fbfcc_buffer <= cw_buffer(49 downto 49);
    -- flow-through slice operator slice_2125_inst
    is_cbccc_buffer <= cw_buffer(48 downto 48);
    -- flow-through slice operator slice_2129_inst
    is_ticc_buffer <= cw_buffer(47 downto 47);
    -- flow-through slice operator slice_2133_inst
    annul_flag_buffer <= cw_buffer(46 downto 46);
    -- flow-through slice operator slice_2137_inst
    br_cond_buffer <= cw_buffer(45 downto 42);
    -- flow-through slice operator slice_2141_inst
    alu_buffer <= cw_buffer(41 downto 41);
    -- flow-through slice operator slice_2145_inst
    use_alu_add_buffer <= cw_buffer(40 downto 40);
    -- flow-through slice operator slice_2149_inst
    is_alu_sub_buffer <= cw_buffer(39 downto 39);
    -- flow-through slice operator slice_2153_inst
    is_alu_mul_buffer <= cw_buffer(38 downto 38);
    -- flow-through slice operator slice_2157_inst
    is_alu_mulscc_buffer <= cw_buffer(37 downto 37);
    -- flow-through slice operator slice_2161_inst
    is_alu_div_buffer <= cw_buffer(36 downto 36);
    -- flow-through slice operator slice_2165_inst
    is_alu_sll_buffer <= cw_buffer(35 downto 35);
    -- flow-through slice operator slice_2169_inst
    is_alu_srl_buffer <= cw_buffer(34 downto 34);
    -- flow-through slice operator slice_2173_inst
    is_alu_sra_buffer <= cw_buffer(33 downto 33);
    -- flow-through slice operator slice_2177_inst
    is_alu_and_buffer <= cw_buffer(32 downto 32);
    -- flow-through slice operator slice_2181_inst
    is_alu_or_buffer <= cw_buffer(31 downto 31);
    -- flow-through slice operator slice_2185_inst
    use_alu_xor_buffer <= cw_buffer(30 downto 30);
    -- flow-through slice operator slice_2189_inst
    is_alu_xnor_buffer <= cw_buffer(29 downto 29);
    -- flow-through slice operator slice_2193_inst
    signed_mul_div_buffer <= cw_buffer(28 downto 28);
    -- flow-through slice operator slice_2197_inst
    negate_second_operand_buffer <= cw_buffer(27 downto 27);
    -- flow-through slice operator slice_2201_inst
    with_carry_buffer <= cw_buffer(26 downto 26);
    -- flow-through slice operator slice_2205_inst
    set_cc_buffer <= cw_buffer(25 downto 25);
    -- flow-through slice operator slice_2209_inst
    tagged_alu_op_buffer <= cw_buffer(24 downto 24);
    -- flow-through slice operator slice_2213_inst
    trap_on_overflow_buffer <= cw_buffer(23 downto 23);
    -- flow-through slice operator slice_2217_inst
    misc_buffer <= cw_buffer(22 downto 22);
    -- flow-through slice operator slice_2221_inst
    is_sethi_buffer <= cw_buffer(21 downto 21);
    -- flow-through slice operator slice_2225_inst
    write_psr_buffer <= cw_buffer(20 downto 20);
    -- flow-through slice operator slice_2229_inst
    write_wim_buffer <= cw_buffer(19 downto 19);
    -- flow-through slice operator slice_2233_inst
    write_tbr_buffer <= cw_buffer(18 downto 18);
    -- flow-through slice operator slice_2237_inst
    write_y_buffer <= cw_buffer(17 downto 17);
    -- flow-through slice operator slice_2241_inst
    write_asr_buffer <= cw_buffer(16 downto 16);
    -- flow-through slice operator slice_2245_inst
    read_psr_buffer <= cw_buffer(15 downto 15);
    -- flow-through slice operator slice_2249_inst
    read_wim_buffer <= cw_buffer(14 downto 14);
    -- flow-through slice operator slice_2253_inst
    read_tbr_buffer <= cw_buffer(13 downto 13);
    -- flow-through slice operator slice_2257_inst
    read_y_buffer <= cw_buffer(12 downto 12);
    -- flow-through slice operator slice_2261_inst
    read_asr_buffer <= cw_buffer(11 downto 11);
    -- flow-through slice operator slice_2265_inst
    asr_id_buffer <= cw_buffer(10 downto 6);
    -- flow-through slice operator slice_2269_inst
    is_save_buffer <= cw_buffer(5 downto 5);
    -- flow-through slice operator slice_2273_inst
    is_restore_buffer <= cw_buffer(4 downto 4);
    -- flow-through slice operator slice_2277_inst
    dti_buffer <= cw_buffer(3 downto 3);
    -- flow-through slice operator slice_2281_inst
    is_iu_dti_buffer <= cw_buffer(2 downto 2);
    -- flow-through slice operator slice_2285_inst
    is_load_to_debug_buffer <= cw_buffer(1 downto 1);
    -- flow-through slice operator slice_2289_inst
    is_store_to_debug_buffer <= cw_buffer(0 downto 0);
    -- 
  end Block; -- data_path
  -- 
end decode_alu_exec_control_word_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity exec_cti_instruction_Volatile is -- 
  port ( -- 
    exec_call : in  std_logic_vector(0 downto 0);
    exec_rett : in  std_logic_vector(0 downto 0);
    exec_jmpl : in  std_logic_vector(0 downto 0);
    exec_ticc : in  std_logic_vector(0 downto 0);
    br_cond : in  std_logic_vector(3 downto 0);
    annul_flag : in  std_logic_vector(0 downto 0);
    pc : in  std_logic_vector(31 downto 0);
    alu_result : in  std_logic_vector(31 downto 0);
    psr : in  std_logic_vector(31 downto 0);
    wim : in  std_logic_vector(31 downto 0);
    cti_trap_status : out  std_logic_vector(0 downto 0);
    cti_ticc_trap_type : out  std_logic_vector(6 downto 0);
    cti_trap_instr_trap : out  std_logic_vector(0 downto 0);
    cti_illegal_instr_trap : out  std_logic_vector(0 downto 0);
    cti_privileged_instr_trap : out  std_logic_vector(0 downto 0);
    cti_window_underflow_trap : out  std_logic_vector(0 downto 0);
    cti_mem_address_not_aligned_trap : out  std_logic_vector(0 downto 0);
    cti_processor_error_mode : out  std_logic_vector(0 downto 0);
    cti_br_taken : out  std_logic_vector(0 downto 0);
    cti_next_psr : out  std_logic_vector(31 downto 0);
    cti_annul_next : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity exec_cti_instruction_Volatile;
architecture exec_cti_instruction_Volatile_arch of exec_cti_instruction_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(137-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal exec_call_buffer :  std_logic_vector(0 downto 0);
  signal exec_rett_buffer :  std_logic_vector(0 downto 0);
  signal exec_jmpl_buffer :  std_logic_vector(0 downto 0);
  signal exec_ticc_buffer :  std_logic_vector(0 downto 0);
  signal br_cond_buffer :  std_logic_vector(3 downto 0);
  signal annul_flag_buffer :  std_logic_vector(0 downto 0);
  signal pc_buffer :  std_logic_vector(31 downto 0);
  signal alu_result_buffer :  std_logic_vector(31 downto 0);
  signal psr_buffer :  std_logic_vector(31 downto 0);
  signal wim_buffer :  std_logic_vector(31 downto 0);
  -- output port buffer signals
  signal cti_trap_status_buffer :  std_logic_vector(0 downto 0);
  signal cti_ticc_trap_type_buffer :  std_logic_vector(6 downto 0);
  signal cti_trap_instr_trap_buffer :  std_logic_vector(0 downto 0);
  signal cti_illegal_instr_trap_buffer :  std_logic_vector(0 downto 0);
  signal cti_privileged_instr_trap_buffer :  std_logic_vector(0 downto 0);
  signal cti_window_underflow_trap_buffer :  std_logic_vector(0 downto 0);
  signal cti_mem_address_not_aligned_trap_buffer :  std_logic_vector(0 downto 0);
  signal cti_processor_error_mode_buffer :  std_logic_vector(0 downto 0);
  signal cti_br_taken_buffer :  std_logic_vector(0 downto 0);
  signal cti_next_psr_buffer :  std_logic_vector(31 downto 0);
  signal cti_annul_next_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  component exec_eval_icc_Volatile is -- 
    port ( -- 
      psr : in  std_logic_vector(31 downto 0);
      br_cond : in  std_logic_vector(3 downto 0);
      annul_flag : in  std_logic_vector(0 downto 0);
      eval_icc : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component exec_rett_instruction_Volatile is -- 
    port ( -- 
      psr : in  std_logic_vector(31 downto 0);
      wim : in  std_logic_vector(31 downto 0);
      alu_result : in  std_logic_vector(31 downto 0);
      new_psr : out  std_logic_vector(31 downto 0);
      rett_trap : out  std_logic_vector(0 downto 0);
      rett_priv_instr_trap : out  std_logic_vector(0 downto 0);
      rett_illegal_instr_trap : out  std_logic_vector(0 downto 0);
      rett_window_underflow_trap : out  std_logic_vector(0 downto 0);
      rett_mem_address_not_aligned_trap : out  std_logic_vector(0 downto 0);
      rett_processor_error_mode : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  exec_call_buffer <= exec_call;
  exec_rett_buffer <= exec_rett;
  exec_jmpl_buffer <= exec_jmpl;
  exec_ticc_buffer <= exec_ticc;
  br_cond_buffer <= br_cond;
  annul_flag_buffer <= annul_flag;
  pc_buffer <= pc;
  alu_result_buffer <= alu_result;
  psr_buffer <= psr;
  wim_buffer <= wim;
  -- output handling  -------------------------------------------------------
  cti_trap_status <= cti_trap_status_buffer;
  cti_ticc_trap_type <= cti_ticc_trap_type_buffer;
  cti_trap_instr_trap <= cti_trap_instr_trap_buffer;
  cti_illegal_instr_trap <= cti_illegal_instr_trap_buffer;
  cti_privileged_instr_trap <= cti_privileged_instr_trap_buffer;
  cti_window_underflow_trap <= cti_window_underflow_trap_buffer;
  cti_mem_address_not_aligned_trap <= cti_mem_address_not_aligned_trap_buffer;
  cti_processor_error_mode <= cti_processor_error_mode_buffer;
  cti_br_taken <= cti_br_taken_buffer;
  cti_next_psr <= cti_next_psr_buffer;
  cti_annul_next <= cti_annul_next_buffer;
  cti_annul_next_buffer <= "0";
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_6490_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6493_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6519_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6544_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6546_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6549_wire : std_logic_vector(0 downto 0);
    signal R_ZERO_7_6510_wire_constant : std_logic_vector(6 downto 0);
    signal eval_icc_6466 : std_logic_vector(0 downto 0);
    signal jmpl_mem_address_not_aligned_trap_6450 : std_logic_vector(0 downto 0);
    signal konst_6448_wire_constant : std_logic_vector(1 downto 0);
    signal new_psr_6461 : std_logic_vector(31 downto 0);
    signal rett_illegal_instr_trap_6461 : std_logic_vector(0 downto 0);
    signal rett_mem_address_not_aligned_trap_6461 : std_logic_vector(0 downto 0);
    signal rett_priv_instr_trap_6461 : std_logic_vector(0 downto 0);
    signal rett_processor_error_mode_6461 : std_logic_vector(0 downto 0);
    signal rett_trap_6461 : std_logic_vector(0 downto 0);
    signal rett_window_underflow_trap_6461 : std_logic_vector(0 downto 0);
    signal slice_6447_wire : std_logic_vector(1 downto 0);
    signal slice_6509_wire : std_logic_vector(6 downto 0);
    signal v_cti_illegal_instr_trap_6476 : std_logic_vector(0 downto 0);
    signal v_cti_mem_address_not_aligned_trap_6495 : std_logic_vector(0 downto 0);
    signal v_cti_privileged_instr_trap_6481 : std_logic_vector(0 downto 0);
    signal v_cti_processor_error_mode_6505 : std_logic_vector(0 downto 0);
    signal v_cti_ticc_trap_instr_trap_6471 : std_logic_vector(0 downto 0);
    signal v_cti_trap_instr_trap_6500 : std_logic_vector(0 downto 0);
    signal v_cti_window_underflow_trap_6486 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_7_6510_wire_constant <= "0000000";
    konst_6448_wire_constant <= "00";
    -- flow-through select operator MUX_6511_inst
    cti_ticc_trap_type_buffer <= slice_6509_wire when (exec_ticc_buffer(0) /=  '0') else R_ZERO_7_6510_wire_constant;
    -- flow-through select operator MUX_6556_inst
    cti_next_psr_buffer <= new_psr_6461 when (exec_rett_buffer(0) /=  '0') else psr_buffer;
    -- flow-through slice operator slice_6447_inst
    slice_6447_wire <= alu_result_buffer(1 downto 0);
    -- flow-through slice operator slice_6509_inst
    slice_6509_wire <= alu_result_buffer(6 downto 0);
    -- interlock W_cti_illegal_instr_trap_6523_inst
    process(v_cti_illegal_instr_trap_6476) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := v_cti_illegal_instr_trap_6476(0 downto 0);
      cti_illegal_instr_trap_buffer <= tmp_var; -- 
    end process;
    -- interlock W_cti_mem_address_not_aligned_trap_6532_inst
    process(v_cti_mem_address_not_aligned_trap_6495) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := v_cti_mem_address_not_aligned_trap_6495(0 downto 0);
      cti_mem_address_not_aligned_trap_buffer <= tmp_var; -- 
    end process;
    -- interlock W_cti_privileged_instr_trap_6526_inst
    process(v_cti_privileged_instr_trap_6481) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := v_cti_privileged_instr_trap_6481(0 downto 0);
      cti_privileged_instr_trap_buffer <= tmp_var; -- 
    end process;
    -- interlock W_cti_processor_error_mode_6538_inst
    process(v_cti_processor_error_mode_6505) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := v_cti_processor_error_mode_6505(0 downto 0);
      cti_processor_error_mode_buffer <= tmp_var; -- 
    end process;
    -- interlock W_cti_trap_instr_trap_6535_inst
    process(v_cti_trap_instr_trap_6500) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := v_cti_trap_instr_trap_6500(0 downto 0);
      cti_trap_instr_trap_buffer <= tmp_var; -- 
    end process;
    -- interlock W_cti_window_underflow_trap_6529_inst
    process(v_cti_window_underflow_trap_6486) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := v_cti_window_underflow_trap_6486(0 downto 0);
      cti_window_underflow_trap_buffer <= tmp_var; -- 
    end process;
    -- flow through binary operator AND_u1_u1_6470_inst
    v_cti_ticc_trap_instr_trap_6471 <= (exec_ticc_buffer and eval_icc_6466);
    -- flow through binary operator AND_u1_u1_6475_inst
    v_cti_illegal_instr_trap_6476 <= (exec_rett_buffer and rett_illegal_instr_trap_6461);
    -- flow through binary operator AND_u1_u1_6480_inst
    v_cti_privileged_instr_trap_6481 <= (exec_rett_buffer and rett_priv_instr_trap_6461);
    -- flow through binary operator AND_u1_u1_6485_inst
    v_cti_window_underflow_trap_6486 <= (exec_rett_buffer and rett_window_underflow_trap_6461);
    -- flow through binary operator AND_u1_u1_6490_inst
    AND_u1_u1_6490_wire <= (exec_rett_buffer and rett_mem_address_not_aligned_trap_6461);
    -- flow through binary operator AND_u1_u1_6493_inst
    AND_u1_u1_6493_wire <= (exec_jmpl_buffer and jmpl_mem_address_not_aligned_trap_6450);
    -- flow through binary operator AND_u1_u1_6499_inst
    v_cti_trap_instr_trap_6500 <= (exec_ticc_buffer and v_cti_ticc_trap_instr_trap_6471);
    -- flow through binary operator AND_u1_u1_6504_inst
    v_cti_processor_error_mode_6505 <= (exec_rett_buffer and rett_processor_error_mode_6461);
    -- flow through binary operator NEQ_u2_u1_6449_inst
    process(slice_6447_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(slice_6447_wire, konst_6448_wire_constant, tmp_var);
      jmpl_mem_address_not_aligned_trap_6450 <= tmp_var; --
    end process;
    -- flow through binary operator OR_u1_u1_6494_inst
    v_cti_mem_address_not_aligned_trap_6495 <= (AND_u1_u1_6490_wire or AND_u1_u1_6493_wire);
    -- flow through binary operator OR_u1_u1_6519_inst
    OR_u1_u1_6519_wire <= (exec_call_buffer or exec_rett_buffer);
    -- flow through binary operator OR_u1_u1_6521_inst
    cti_br_taken_buffer <= (OR_u1_u1_6519_wire or exec_jmpl_buffer);
    -- flow through binary operator OR_u1_u1_6544_inst
    OR_u1_u1_6544_wire <= (v_cti_illegal_instr_trap_6476 or v_cti_privileged_instr_trap_6481);
    -- flow through binary operator OR_u1_u1_6546_inst
    OR_u1_u1_6546_wire <= (OR_u1_u1_6544_wire or v_cti_window_underflow_trap_6486);
    -- flow through binary operator OR_u1_u1_6549_inst
    OR_u1_u1_6549_wire <= (v_cti_mem_address_not_aligned_trap_6495 or v_cti_trap_instr_trap_6500);
    -- flow through binary operator OR_u1_u1_6550_inst
    cti_trap_status_buffer <= (OR_u1_u1_6546_wire or OR_u1_u1_6549_wire);
    volatile_operator_exec_rett_instruction_5390: exec_rett_instruction_Volatile port map(psr => psr_buffer, wim => wim_buffer, alu_result => alu_result_buffer, new_psr => new_psr_6461, rett_trap => rett_trap_6461, rett_priv_instr_trap => rett_priv_instr_trap_6461, rett_illegal_instr_trap => rett_illegal_instr_trap_6461, rett_window_underflow_trap => rett_window_underflow_trap_6461, rett_mem_address_not_aligned_trap => rett_mem_address_not_aligned_trap_6461, rett_processor_error_mode => rett_processor_error_mode_6461); 
    volatile_operator_exec_eval_icc_5391: exec_eval_icc_Volatile port map(psr => psr_buffer, br_cond => br_cond_buffer, annul_flag => annul_flag_buffer, eval_icc => eval_icc_6466); 
    -- 
  end Block; -- data_path
  -- 
end exec_cti_instruction_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity exec_eval_icc_Volatile is -- 
  port ( -- 
    psr : in  std_logic_vector(31 downto 0);
    br_cond : in  std_logic_vector(3 downto 0);
    annul_flag : in  std_logic_vector(0 downto 0);
    eval_icc : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity exec_eval_icc_Volatile;
architecture exec_eval_icc_Volatile_arch of exec_eval_icc_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(37-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal psr_buffer :  std_logic_vector(31 downto 0);
  signal br_cond_buffer :  std_logic_vector(3 downto 0);
  signal annul_flag_buffer :  std_logic_vector(0 downto 0);
  -- output port buffer signals
  signal eval_icc_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  psr_buffer <= psr;
  br_cond_buffer <= br_cond;
  annul_flag_buffer <= annul_flag;
  -- output handling  -------------------------------------------------------
  eval_icc <= eval_icc_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal C_6285 : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6289_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6295_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6302_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6309_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6317_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6328_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6339_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6348_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6359_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6368_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6377_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6384_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6392_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6399_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6406_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_6413_wire : std_logic_vector(0 downto 0);
    signal MUX_6292_wire : std_logic_vector(0 downto 0);
    signal MUX_6298_wire : std_logic_vector(0 downto 0);
    signal MUX_6306_wire : std_logic_vector(0 downto 0);
    signal MUX_6312_wire : std_logic_vector(0 downto 0);
    signal MUX_6325_wire : std_logic_vector(0 downto 0);
    signal MUX_6335_wire : std_logic_vector(0 downto 0);
    signal MUX_6345_wire : std_logic_vector(0 downto 0);
    signal MUX_6353_wire : std_logic_vector(0 downto 0);
    signal MUX_6365_wire : std_logic_vector(0 downto 0);
    signal MUX_6373_wire : std_logic_vector(0 downto 0);
    signal MUX_6381_wire : std_logic_vector(0 downto 0);
    signal MUX_6387_wire : std_logic_vector(0 downto 0);
    signal MUX_6396_wire : std_logic_vector(0 downto 0);
    signal MUX_6402_wire : std_logic_vector(0 downto 0);
    signal MUX_6410_wire : std_logic_vector(0 downto 0);
    signal MUX_6416_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6304_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6323_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6343_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6363_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6379_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6394_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6408_wire : std_logic_vector(0 downto 0);
    signal N_6270 : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6299_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6313_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6314_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6322_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6333_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6336_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6354_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6355_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6356_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6362_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6371_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6374_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6388_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6389_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6403_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6417_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6418_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6419_wire : std_logic_vector(0 downto 0);
    signal R_ONE_1_6290_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_6296_wire_constant : std_logic_vector(0 downto 0);
    signal V_6280 : std_logic_vector(0 downto 0);
    signal XOR_u1_u1_6321_wire : std_logic_vector(0 downto 0);
    signal XOR_u1_u1_6332_wire : std_logic_vector(0 downto 0);
    signal XOR_u1_u1_6342_wire : std_logic_vector(0 downto 0);
    signal XOR_u1_u1_6351_wire : std_logic_vector(0 downto 0);
    signal Z_6275 : std_logic_vector(0 downto 0);
    signal konst_6268_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6273_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6278_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6283_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6288_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6291_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6294_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6297_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6301_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6305_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6308_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6311_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6316_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6324_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6327_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6334_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6338_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6344_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6347_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6352_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6358_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6364_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6367_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6372_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6376_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6380_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6383_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6386_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6391_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6395_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6398_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6401_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6405_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6409_wire_constant : std_logic_vector(0 downto 0);
    signal konst_6412_wire_constant : std_logic_vector(3 downto 0);
    signal konst_6415_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ONE_1_6290_wire_constant <= "1";
    R_ZERO_1_6296_wire_constant <= "0";
    konst_6268_wire_constant <= "00000000000000000000000000010111";
    konst_6273_wire_constant <= "00000000000000000000000000010110";
    konst_6278_wire_constant <= "00000000000000000000000000010101";
    konst_6283_wire_constant <= "00000000000000000000000000010100";
    konst_6288_wire_constant <= "1000";
    konst_6291_wire_constant <= "0";
    konst_6294_wire_constant <= "0000";
    konst_6297_wire_constant <= "0";
    konst_6301_wire_constant <= "1001";
    konst_6305_wire_constant <= "0";
    konst_6308_wire_constant <= "0001";
    konst_6311_wire_constant <= "0";
    konst_6316_wire_constant <= "1010";
    konst_6324_wire_constant <= "0";
    konst_6327_wire_constant <= "0010";
    konst_6334_wire_constant <= "0";
    konst_6338_wire_constant <= "1011";
    konst_6344_wire_constant <= "0";
    konst_6347_wire_constant <= "0011";
    konst_6352_wire_constant <= "0";
    konst_6358_wire_constant <= "1100";
    konst_6364_wire_constant <= "0";
    konst_6367_wire_constant <= "0100";
    konst_6372_wire_constant <= "0";
    konst_6376_wire_constant <= "1101";
    konst_6380_wire_constant <= "0";
    konst_6383_wire_constant <= "0101";
    konst_6386_wire_constant <= "0";
    konst_6391_wire_constant <= "1110";
    konst_6395_wire_constant <= "0";
    konst_6398_wire_constant <= "0110";
    konst_6401_wire_constant <= "0";
    konst_6405_wire_constant <= "1111";
    konst_6409_wire_constant <= "0";
    konst_6412_wire_constant <= "0111";
    konst_6415_wire_constant <= "0";
    -- flow-through select operator MUX_6292_inst
    MUX_6292_wire <= R_ONE_1_6290_wire_constant when (EQ_u4_u1_6289_wire(0) /=  '0') else konst_6291_wire_constant;
    -- flow-through select operator MUX_6298_inst
    MUX_6298_wire <= R_ZERO_1_6296_wire_constant when (EQ_u4_u1_6295_wire(0) /=  '0') else konst_6297_wire_constant;
    -- flow-through select operator MUX_6306_inst
    MUX_6306_wire <= NOT_u1_u1_6304_wire when (EQ_u4_u1_6302_wire(0) /=  '0') else konst_6305_wire_constant;
    -- flow-through select operator MUX_6312_inst
    MUX_6312_wire <= Z_6275 when (EQ_u4_u1_6309_wire(0) /=  '0') else konst_6311_wire_constant;
    -- flow-through select operator MUX_6325_inst
    MUX_6325_wire <= NOT_u1_u1_6323_wire when (EQ_u4_u1_6317_wire(0) /=  '0') else konst_6324_wire_constant;
    -- flow-through select operator MUX_6335_inst
    MUX_6335_wire <= OR_u1_u1_6333_wire when (EQ_u4_u1_6328_wire(0) /=  '0') else konst_6334_wire_constant;
    -- flow-through select operator MUX_6345_inst
    MUX_6345_wire <= NOT_u1_u1_6343_wire when (EQ_u4_u1_6339_wire(0) /=  '0') else konst_6344_wire_constant;
    -- flow-through select operator MUX_6353_inst
    MUX_6353_wire <= XOR_u1_u1_6351_wire when (EQ_u4_u1_6348_wire(0) /=  '0') else konst_6352_wire_constant;
    -- flow-through select operator MUX_6365_inst
    MUX_6365_wire <= NOT_u1_u1_6363_wire when (EQ_u4_u1_6359_wire(0) /=  '0') else konst_6364_wire_constant;
    -- flow-through select operator MUX_6373_inst
    MUX_6373_wire <= OR_u1_u1_6371_wire when (EQ_u4_u1_6368_wire(0) /=  '0') else konst_6372_wire_constant;
    -- flow-through select operator MUX_6381_inst
    MUX_6381_wire <= NOT_u1_u1_6379_wire when (EQ_u4_u1_6377_wire(0) /=  '0') else konst_6380_wire_constant;
    -- flow-through select operator MUX_6387_inst
    MUX_6387_wire <= C_6285 when (EQ_u4_u1_6384_wire(0) /=  '0') else konst_6386_wire_constant;
    -- flow-through select operator MUX_6396_inst
    MUX_6396_wire <= NOT_u1_u1_6394_wire when (EQ_u4_u1_6392_wire(0) /=  '0') else konst_6395_wire_constant;
    -- flow-through select operator MUX_6402_inst
    MUX_6402_wire <= N_6270 when (EQ_u4_u1_6399_wire(0) /=  '0') else konst_6401_wire_constant;
    -- flow-through select operator MUX_6410_inst
    MUX_6410_wire <= NOT_u1_u1_6408_wire when (EQ_u4_u1_6406_wire(0) /=  '0') else konst_6409_wire_constant;
    -- flow-through select operator MUX_6416_inst
    MUX_6416_wire <= V_6280 when (EQ_u4_u1_6413_wire(0) /=  '0') else konst_6415_wire_constant;
    -- flow through binary operator BITSEL_u32_u1_6269_inst
    process(psr_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(psr_buffer, konst_6268_wire_constant, tmp_var);
      N_6270 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6274_inst
    process(psr_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(psr_buffer, konst_6273_wire_constant, tmp_var);
      Z_6275 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6279_inst
    process(psr_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(psr_buffer, konst_6278_wire_constant, tmp_var);
      V_6280 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6284_inst
    process(psr_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(psr_buffer, konst_6283_wire_constant, tmp_var);
      C_6285 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6289_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6288_wire_constant, tmp_var);
      EQ_u4_u1_6289_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6295_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6294_wire_constant, tmp_var);
      EQ_u4_u1_6295_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6302_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6301_wire_constant, tmp_var);
      EQ_u4_u1_6302_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6309_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6308_wire_constant, tmp_var);
      EQ_u4_u1_6309_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6317_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6316_wire_constant, tmp_var);
      EQ_u4_u1_6317_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6328_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6327_wire_constant, tmp_var);
      EQ_u4_u1_6328_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6339_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6338_wire_constant, tmp_var);
      EQ_u4_u1_6339_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6348_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6347_wire_constant, tmp_var);
      EQ_u4_u1_6348_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6359_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6358_wire_constant, tmp_var);
      EQ_u4_u1_6359_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6368_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6367_wire_constant, tmp_var);
      EQ_u4_u1_6368_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6377_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6376_wire_constant, tmp_var);
      EQ_u4_u1_6377_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6384_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6383_wire_constant, tmp_var);
      EQ_u4_u1_6384_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6392_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6391_wire_constant, tmp_var);
      EQ_u4_u1_6392_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6399_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6398_wire_constant, tmp_var);
      EQ_u4_u1_6399_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6406_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6405_wire_constant, tmp_var);
      EQ_u4_u1_6406_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_6413_inst
    process(br_cond_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(br_cond_buffer, konst_6412_wire_constant, tmp_var);
      EQ_u4_u1_6413_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_6304_inst
    process(Z_6275) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", Z_6275, tmp_var);
      NOT_u1_u1_6304_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6323_inst
    process(OR_u1_u1_6322_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", OR_u1_u1_6322_wire, tmp_var);
      NOT_u1_u1_6323_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6343_inst
    process(XOR_u1_u1_6342_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", XOR_u1_u1_6342_wire, tmp_var);
      NOT_u1_u1_6343_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6363_inst
    process(OR_u1_u1_6362_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", OR_u1_u1_6362_wire, tmp_var);
      NOT_u1_u1_6363_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6379_inst
    process(C_6285) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", C_6285, tmp_var);
      NOT_u1_u1_6379_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6394_inst
    process(N_6270) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", N_6270, tmp_var);
      NOT_u1_u1_6394_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6408_inst
    process(V_6280) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", V_6280, tmp_var);
      NOT_u1_u1_6408_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_6299_inst
    OR_u1_u1_6299_wire <= (MUX_6292_wire or MUX_6298_wire);
    -- flow through binary operator OR_u1_u1_6313_inst
    OR_u1_u1_6313_wire <= (MUX_6306_wire or MUX_6312_wire);
    -- flow through binary operator OR_u1_u1_6314_inst
    OR_u1_u1_6314_wire <= (OR_u1_u1_6299_wire or OR_u1_u1_6313_wire);
    -- flow through binary operator OR_u1_u1_6322_inst
    OR_u1_u1_6322_wire <= (Z_6275 or XOR_u1_u1_6321_wire);
    -- flow through binary operator OR_u1_u1_6333_inst
    OR_u1_u1_6333_wire <= (Z_6275 or XOR_u1_u1_6332_wire);
    -- flow through binary operator OR_u1_u1_6336_inst
    OR_u1_u1_6336_wire <= (MUX_6325_wire or MUX_6335_wire);
    -- flow through binary operator OR_u1_u1_6354_inst
    OR_u1_u1_6354_wire <= (MUX_6345_wire or MUX_6353_wire);
    -- flow through binary operator OR_u1_u1_6355_inst
    OR_u1_u1_6355_wire <= (OR_u1_u1_6336_wire or OR_u1_u1_6354_wire);
    -- flow through binary operator OR_u1_u1_6356_inst
    OR_u1_u1_6356_wire <= (OR_u1_u1_6314_wire or OR_u1_u1_6355_wire);
    -- flow through binary operator OR_u1_u1_6362_inst
    OR_u1_u1_6362_wire <= (C_6285 or Z_6275);
    -- flow through binary operator OR_u1_u1_6371_inst
    OR_u1_u1_6371_wire <= (C_6285 or Z_6275);
    -- flow through binary operator OR_u1_u1_6374_inst
    OR_u1_u1_6374_wire <= (MUX_6365_wire or MUX_6373_wire);
    -- flow through binary operator OR_u1_u1_6388_inst
    OR_u1_u1_6388_wire <= (MUX_6381_wire or MUX_6387_wire);
    -- flow through binary operator OR_u1_u1_6389_inst
    OR_u1_u1_6389_wire <= (OR_u1_u1_6374_wire or OR_u1_u1_6388_wire);
    -- flow through binary operator OR_u1_u1_6403_inst
    OR_u1_u1_6403_wire <= (MUX_6396_wire or MUX_6402_wire);
    -- flow through binary operator OR_u1_u1_6417_inst
    OR_u1_u1_6417_wire <= (MUX_6410_wire or MUX_6416_wire);
    -- flow through binary operator OR_u1_u1_6418_inst
    OR_u1_u1_6418_wire <= (OR_u1_u1_6403_wire or OR_u1_u1_6417_wire);
    -- flow through binary operator OR_u1_u1_6419_inst
    OR_u1_u1_6419_wire <= (OR_u1_u1_6389_wire or OR_u1_u1_6418_wire);
    -- flow through binary operator OR_u1_u1_6420_inst
    eval_icc_buffer <= (OR_u1_u1_6356_wire or OR_u1_u1_6419_wire);
    -- flow through binary operator XOR_u1_u1_6321_inst
    XOR_u1_u1_6321_wire <= (N_6270 xor V_6280);
    -- flow through binary operator XOR_u1_u1_6332_inst
    XOR_u1_u1_6332_wire <= (N_6270 xor V_6280);
    -- flow through binary operator XOR_u1_u1_6342_inst
    XOR_u1_u1_6342_wire <= (N_6270 xor V_6280);
    -- flow through binary operator XOR_u1_u1_6351_inst
    XOR_u1_u1_6351_wire <= (N_6270 xor V_6280);
    -- 
  end Block; -- data_path
  -- 
end exec_eval_icc_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity exec_rett_instruction_Volatile is -- 
  port ( -- 
    psr : in  std_logic_vector(31 downto 0);
    wim : in  std_logic_vector(31 downto 0);
    alu_result : in  std_logic_vector(31 downto 0);
    new_psr : out  std_logic_vector(31 downto 0);
    rett_trap : out  std_logic_vector(0 downto 0);
    rett_priv_instr_trap : out  std_logic_vector(0 downto 0);
    rett_illegal_instr_trap : out  std_logic_vector(0 downto 0);
    rett_window_underflow_trap : out  std_logic_vector(0 downto 0);
    rett_mem_address_not_aligned_trap : out  std_logic_vector(0 downto 0);
    rett_processor_error_mode : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity exec_rett_instruction_Volatile;
architecture exec_rett_instruction_Volatile_arch of exec_rett_instruction_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(96-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal psr_buffer :  std_logic_vector(31 downto 0);
  signal wim_buffer :  std_logic_vector(31 downto 0);
  signal alu_result_buffer :  std_logic_vector(31 downto 0);
  -- output port buffer signals
  signal new_psr_buffer :  std_logic_vector(31 downto 0);
  signal rett_trap_buffer :  std_logic_vector(0 downto 0);
  signal rett_priv_instr_trap_buffer :  std_logic_vector(0 downto 0);
  signal rett_illegal_instr_trap_buffer :  std_logic_vector(0 downto 0);
  signal rett_window_underflow_trap_buffer :  std_logic_vector(0 downto 0);
  signal rett_mem_address_not_aligned_trap_buffer :  std_logic_vector(0 downto 0);
  signal rett_processor_error_mode_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  psr_buffer <= psr;
  wim_buffer <= wim;
  alu_result_buffer <= alu_result;
  -- output handling  -------------------------------------------------------
  new_psr <= new_psr_buffer;
  rett_trap <= rett_trap_buffer;
  rett_priv_instr_trap <= rett_priv_instr_trap_buffer;
  rett_illegal_instr_trap <= rett_illegal_instr_trap_buffer;
  rett_window_underflow_trap <= rett_window_underflow_trap_buffer;
  rett_mem_address_not_aligned_trap <= rett_mem_address_not_aligned_trap_buffer;
  rett_processor_error_mode <= rett_processor_error_mode_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal ADD_u5_u5_6123_wire : std_logic_vector(4 downto 0);
    signal AND_u32_u32_6167_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u1_u6_6245_wire : std_logic_vector(5 downto 0);
    signal CONCAT_u24_u25_6240_wire : std_logic_vector(24 downto 0);
    signal CONCAT_u25_u26_6242_wire : std_logic_vector(25 downto 0);
    signal MUX_6153_wire : std_logic_vector(0 downto 0);
    signal MUX_6180_wire : std_logic_vector(0 downto 0);
    signal MUX_6181_wire : std_logic_vector(0 downto 0);
    signal MUX_6198_wire : std_logic_vector(0 downto 0);
    signal MUX_6199_wire : std_logic_vector(0 downto 0);
    signal MUX_6200_wire : std_logic_vector(0 downto 0);
    signal MUX_6217_wire : std_logic_vector(0 downto 0);
    signal MUX_6218_wire : std_logic_vector(0 downto 0);
    signal MUX_6219_wire : std_logic_vector(0 downto 0);
    signal NEQ_u2_u1_6195_wire : std_logic_vector(0 downto 0);
    signal NEQ_u2_u1_6214_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6148_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6150_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6175_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6188_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6207_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6225_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6227_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6230_wire : std_logic_vector(0 downto 0);
    signal PS_6141 : std_logic_vector(0 downto 0);
    signal R_NWINDOWS_MOD_MASK_5_6124_wire_constant : std_logic_vector(4 downto 0);
    signal R_ONE_1_6151_wire_constant : std_logic_vector(0 downto 0);
    signal R_ONE_1_6178_wire_constant : std_logic_vector(0 downto 0);
    signal R_ONE_1_6196_wire_constant : std_logic_vector(0 downto 0);
    signal R_ONE_1_6208_wire_constant : std_logic_vector(0 downto 0);
    signal R_ONE_1_6210_wire_constant : std_logic_vector(0 downto 0);
    signal R_ONE_1_6215_wire_constant : std_logic_vector(0 downto 0);
    signal R_ONE_32_6163_wire_constant : std_logic_vector(31 downto 0);
    signal R_ZERO_1_6152_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_6173_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_6176_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_6179_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_6186_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_6189_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_6191_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_6197_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_6205_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_6216_wire_constant : std_logic_vector(0 downto 0);
    signal SHL_u32_u32_6166_wire : std_logic_vector(31 downto 0);
    signal S_6136 : std_logic_vector(0 downto 0);
    signal cwp_6119 : std_logic_vector(4 downto 0);
    signal et_6131 : std_logic_vector(0 downto 0);
    signal konst_6122_wire_constant : std_logic_vector(4 downto 0);
    signal konst_6129_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6134_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6139_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6168_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6194_wire_constant : std_logic_vector(1 downto 0);
    signal konst_6213_wire_constant : std_logic_vector(1 downto 0);
    signal nET_6235 : std_logic_vector(0 downto 0);
    signal nS_6144 : std_logic_vector(0 downto 0);
    signal new_cwp_6126 : std_logic_vector(4 downto 0);
    signal slice_6193_wire : std_logic_vector(1 downto 0);
    signal slice_6212_wire : std_logic_vector(1 downto 0);
    signal slice_6238_wire : std_logic_vector(23 downto 0);
    signal type_cast_6165_wire : std_logic_vector(31 downto 0);
    signal wim_cwp_flag_6170 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_NWINDOWS_MOD_MASK_5_6124_wire_constant <= "00111";
    R_ONE_1_6151_wire_constant <= "1";
    R_ONE_1_6178_wire_constant <= "1";
    R_ONE_1_6196_wire_constant <= "1";
    R_ONE_1_6208_wire_constant <= "1";
    R_ONE_1_6210_wire_constant <= "1";
    R_ONE_1_6215_wire_constant <= "1";
    R_ONE_32_6163_wire_constant <= "00000000000000000000000000000001";
    R_ZERO_1_6152_wire_constant <= "0";
    R_ZERO_1_6173_wire_constant <= "0";
    R_ZERO_1_6176_wire_constant <= "0";
    R_ZERO_1_6179_wire_constant <= "0";
    R_ZERO_1_6186_wire_constant <= "0";
    R_ZERO_1_6189_wire_constant <= "0";
    R_ZERO_1_6191_wire_constant <= "0";
    R_ZERO_1_6197_wire_constant <= "0";
    R_ZERO_1_6205_wire_constant <= "0";
    R_ZERO_1_6216_wire_constant <= "0";
    konst_6122_wire_constant <= "00001";
    konst_6129_wire_constant <= "00000000000000000000000000000101";
    konst_6134_wire_constant <= "00000000000000000000000000000111";
    konst_6139_wire_constant <= "00000000000000000000000000000110";
    konst_6168_wire_constant <= "00000000000000000000000000000000";
    konst_6194_wire_constant <= "00";
    konst_6213_wire_constant <= "00";
    nET_6235 <= "1";
    -- flow-through select operator MUX_6153_inst
    MUX_6153_wire <= R_ONE_1_6151_wire_constant when (NOT_u1_u1_6150_wire(0) /=  '0') else R_ZERO_1_6152_wire_constant;
    -- flow-through select operator MUX_6154_inst
    rett_priv_instr_trap_buffer <= NOT_u1_u1_6148_wire when (et_6131(0) /=  '0') else MUX_6153_wire;
    -- flow-through select operator MUX_6180_inst
    MUX_6180_wire <= R_ONE_1_6178_wire_constant when (wim_cwp_flag_6170(0) /=  '0') else R_ZERO_1_6179_wire_constant;
    -- flow-through select operator MUX_6181_inst
    MUX_6181_wire <= R_ZERO_1_6176_wire_constant when (NOT_u1_u1_6175_wire(0) /=  '0') else MUX_6180_wire;
    -- flow-through select operator MUX_6182_inst
    rett_window_underflow_trap_buffer <= R_ZERO_1_6173_wire_constant when (et_6131(0) /=  '0') else MUX_6181_wire;
    -- flow-through select operator MUX_6198_inst
    MUX_6198_wire <= R_ONE_1_6196_wire_constant when (NEQ_u2_u1_6195_wire(0) /=  '0') else R_ZERO_1_6197_wire_constant;
    -- flow-through select operator MUX_6199_inst
    MUX_6199_wire <= R_ZERO_1_6191_wire_constant when (wim_cwp_flag_6170(0) /=  '0') else MUX_6198_wire;
    -- flow-through select operator MUX_6200_inst
    MUX_6200_wire <= R_ZERO_1_6189_wire_constant when (NOT_u1_u1_6188_wire(0) /=  '0') else MUX_6199_wire;
    -- flow-through select operator MUX_6201_inst
    rett_mem_address_not_aligned_trap_buffer <= R_ZERO_1_6186_wire_constant when (et_6131(0) /=  '0') else MUX_6200_wire;
    -- flow-through select operator MUX_6217_inst
    MUX_6217_wire <= R_ONE_1_6215_wire_constant when (NEQ_u2_u1_6214_wire(0) /=  '0') else R_ZERO_1_6216_wire_constant;
    -- flow-through select operator MUX_6218_inst
    MUX_6218_wire <= R_ONE_1_6210_wire_constant when (wim_cwp_flag_6170(0) /=  '0') else MUX_6217_wire;
    -- flow-through select operator MUX_6219_inst
    MUX_6219_wire <= R_ONE_1_6208_wire_constant when (NOT_u1_u1_6207_wire(0) /=  '0') else MUX_6218_wire;
    -- flow-through select operator MUX_6220_inst
    rett_processor_error_mode_buffer <= R_ZERO_1_6205_wire_constant when (et_6131(0) /=  '0') else MUX_6219_wire;
    -- flow-through slice operator slice_6118_inst
    cwp_6119 <= psr_buffer(4 downto 0);
    -- flow-through slice operator slice_6193_inst
    slice_6193_wire <= alu_result_buffer(1 downto 0);
    -- flow-through slice operator slice_6212_inst
    slice_6212_wire <= alu_result_buffer(1 downto 0);
    -- flow-through slice operator slice_6238_inst
    slice_6238_wire <= psr_buffer(31 downto 8);
    -- interlock W_nS_6142_inst
    process(PS_6141) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := PS_6141(0 downto 0);
      nS_6144 <= tmp_var; -- 
    end process;
    -- interlock type_cast_6165_inst
    process(new_cwp_6126) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 4 downto 0) := new_cwp_6126(4 downto 0);
      type_cast_6165_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator ADD_u5_u5_6123_inst
    ADD_u5_u5_6123_wire <= std_logic_vector(unsigned(cwp_6119) + unsigned(konst_6122_wire_constant));
    -- flow through binary operator AND_u1_u1_6159_inst
    rett_illegal_instr_trap_buffer <= (et_6131 and S_6136);
    -- flow through binary operator AND_u32_u32_6167_inst
    AND_u32_u32_6167_wire <= (wim_buffer and SHL_u32_u32_6166_wire);
    -- flow through binary operator AND_u5_u5_6125_inst
    new_cwp_6126 <= (ADD_u5_u5_6123_wire and R_NWINDOWS_MOD_MASK_5_6124_wire_constant);
    -- flow through binary operator BITSEL_u32_u1_6130_inst
    process(psr_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(psr_buffer, konst_6129_wire_constant, tmp_var);
      et_6131 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6135_inst
    process(psr_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(psr_buffer, konst_6134_wire_constant, tmp_var);
      S_6136 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6140_inst
    process(psr_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(psr_buffer, konst_6139_wire_constant, tmp_var);
      PS_6141 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u6_6245_inst
    process(nET_6235, new_cwp_6126) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(nET_6235, new_cwp_6126, tmp_var);
      CONCAT_u1_u6_6245_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u24_u25_6240_inst
    process(slice_6238_wire, nS_6144) -- 
      variable tmp_var : std_logic_vector(24 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_6238_wire, nS_6144, tmp_var);
      CONCAT_u24_u25_6240_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u25_u26_6242_inst
    process(CONCAT_u24_u25_6240_wire, PS_6141) -- 
      variable tmp_var : std_logic_vector(25 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u24_u25_6240_wire, PS_6141, tmp_var);
      CONCAT_u25_u26_6242_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u26_u32_6246_inst
    process(CONCAT_u25_u26_6242_wire, CONCAT_u1_u6_6245_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u25_u26_6242_wire, CONCAT_u1_u6_6245_wire, tmp_var);
      new_psr_buffer <= tmp_var; --
    end process;
    -- flow through binary operator NEQ_u2_u1_6195_inst
    process(slice_6193_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(slice_6193_wire, konst_6194_wire_constant, tmp_var);
      NEQ_u2_u1_6195_wire <= tmp_var; --
    end process;
    -- flow through binary operator NEQ_u2_u1_6214_inst
    process(slice_6212_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(slice_6212_wire, konst_6213_wire_constant, tmp_var);
      NEQ_u2_u1_6214_wire <= tmp_var; --
    end process;
    -- flow through binary operator NEQ_u32_u1_6169_inst
    process(AND_u32_u32_6167_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(AND_u32_u32_6167_wire, konst_6168_wire_constant, tmp_var);
      wim_cwp_flag_6170 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_6148_inst
    process(S_6136) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", S_6136, tmp_var);
      NOT_u1_u1_6148_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6150_inst
    process(S_6136) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", S_6136, tmp_var);
      NOT_u1_u1_6150_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6175_inst
    process(S_6136) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", S_6136, tmp_var);
      NOT_u1_u1_6175_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6188_inst
    process(S_6136) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", S_6136, tmp_var);
      NOT_u1_u1_6188_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6207_inst
    process(S_6136) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", S_6136, tmp_var);
      NOT_u1_u1_6207_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_6225_inst
    OR_u1_u1_6225_wire <= (rett_priv_instr_trap_buffer or rett_illegal_instr_trap_buffer);
    -- flow through binary operator OR_u1_u1_6227_inst
    OR_u1_u1_6227_wire <= (OR_u1_u1_6225_wire or rett_window_underflow_trap_buffer);
    -- flow through binary operator OR_u1_u1_6230_inst
    OR_u1_u1_6230_wire <= (rett_mem_address_not_aligned_trap_buffer or rett_processor_error_mode_buffer);
    -- flow through binary operator OR_u1_u1_6231_inst
    rett_trap_buffer <= (OR_u1_u1_6227_wire or OR_u1_u1_6230_wire);
    -- flow through binary operator SHL_u32_u32_6166_inst
    process(R_ONE_32_6163_wire_constant, type_cast_6165_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(R_ONE_32_6163_wire_constant, type_cast_6165_wire, tmp_var);
      SHL_u32_u32_6166_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end exec_rett_instruction_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity find_left_16_Volatile is -- 
  port ( -- 
    fp_16 : in  std_logic_vector(15 downto 0);
    position : out  std_logic_vector(3 downto 0);
    found : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity find_left_16_Volatile;
architecture find_left_16_Volatile_arch of find_left_16_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(16-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal fp_16_buffer :  std_logic_vector(15 downto 0);
  -- output port buffer signals
  signal position_buffer :  std_logic_vector(3 downto 0);
  signal found_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  component find_left_8_Volatile is -- 
    port ( -- 
      fp_8 : in  std_logic_vector(7 downto 0);
      position : out  std_logic_vector(2 downto 0);
      found : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  fp_16_buffer <= fp_16;
  -- output handling  -------------------------------------------------------
  position <= position_buffer;
  found <= found_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u4_1105_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u1_u4_1109_wire : std_logic_vector(3 downto 0);
    signal MUX_1111_wire : std_logic_vector(3 downto 0);
    signal R_ONE_1_1103_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_1107_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_4_1110_wire_constant : std_logic_vector(3 downto 0);
    signal found_lower_1100 : std_logic_vector(0 downto 0);
    signal found_upper_1096 : std_logic_vector(0 downto 0);
    signal fp_8_lower_1092 : std_logic_vector(7 downto 0);
    signal fp_8_lower_index_1100 : std_logic_vector(2 downto 0);
    signal fp_8_upper_1088 : std_logic_vector(7 downto 0);
    signal fp_8_upper_index_1096 : std_logic_vector(2 downto 0);
    -- 
  begin -- 
    R_ONE_1_1103_wire_constant <= "1";
    R_ZERO_1_1107_wire_constant <= "0";
    R_ZERO_4_1110_wire_constant <= "0000";
    -- flow-through select operator MUX_1111_inst
    MUX_1111_wire <= CONCAT_u1_u4_1109_wire when (found_lower_1100(0) /=  '0') else R_ZERO_4_1110_wire_constant;
    -- flow-through select operator MUX_1112_inst
    position_buffer <= CONCAT_u1_u4_1105_wire when (found_upper_1096(0) /=  '0') else MUX_1111_wire;
    -- flow-through slice operator slice_1087_inst
    fp_8_upper_1088 <= fp_16_buffer(15 downto 8);
    -- flow-through slice operator slice_1091_inst
    fp_8_lower_1092 <= fp_16_buffer(7 downto 0);
    -- flow through binary operator CONCAT_u1_u4_1105_inst
    process(R_ONE_1_1103_wire_constant, fp_8_upper_index_1096) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_1103_wire_constant, fp_8_upper_index_1096, tmp_var);
      CONCAT_u1_u4_1105_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u4_1109_inst
    process(R_ZERO_1_1107_wire_constant, fp_8_lower_index_1100) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_1_1107_wire_constant, fp_8_lower_index_1100, tmp_var);
      CONCAT_u1_u4_1109_wire <= tmp_var; --
    end process;
    -- flow through binary operator OR_u1_u1_1117_inst
    found_buffer <= (found_upper_1096 or found_lower_1100);
    volatile_operator_find_left_8_767: find_left_8_Volatile port map(fp_8 => fp_8_upper_1088, position => fp_8_upper_index_1096, found => found_upper_1096); 
    volatile_operator_find_left_8_768: find_left_8_Volatile port map(fp_8 => fp_8_lower_1092, position => fp_8_lower_index_1100, found => found_lower_1100); 
    -- 
  end Block; -- data_path
  -- 
end find_left_16_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity find_left_32_Volatile is -- 
  port ( -- 
    fp_32 : in  std_logic_vector(31 downto 0);
    position : out  std_logic_vector(4 downto 0);
    found : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity find_left_32_Volatile;
architecture find_left_32_Volatile_arch of find_left_32_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(32-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal fp_32_buffer :  std_logic_vector(31 downto 0);
  -- output port buffer signals
  signal position_buffer :  std_logic_vector(4 downto 0);
  signal found_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  component find_left_16_Volatile is -- 
    port ( -- 
      fp_16 : in  std_logic_vector(15 downto 0);
      position : out  std_logic_vector(3 downto 0);
      found : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  fp_32_buffer <= fp_32;
  -- output handling  -------------------------------------------------------
  position <= position_buffer;
  found <= found_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u5_1144_wire : std_logic_vector(4 downto 0);
    signal CONCAT_u1_u5_1148_wire : std_logic_vector(4 downto 0);
    signal MUX_1150_wire : std_logic_vector(4 downto 0);
    signal R_ONE_1_1142_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_1146_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_5_1149_wire_constant : std_logic_vector(4 downto 0);
    signal found_lower_1139 : std_logic_vector(0 downto 0);
    signal found_upper_1135 : std_logic_vector(0 downto 0);
    signal fp_16_lower_1131 : std_logic_vector(15 downto 0);
    signal fp_16_lower_index_1139 : std_logic_vector(3 downto 0);
    signal fp_16_upper_1127 : std_logic_vector(15 downto 0);
    signal fp_16_upper_index_1135 : std_logic_vector(3 downto 0);
    -- 
  begin -- 
    R_ONE_1_1142_wire_constant <= "1";
    R_ZERO_1_1146_wire_constant <= "0";
    R_ZERO_5_1149_wire_constant <= "00000";
    -- flow-through select operator MUX_1150_inst
    MUX_1150_wire <= CONCAT_u1_u5_1148_wire when (found_lower_1139(0) /=  '0') else R_ZERO_5_1149_wire_constant;
    -- flow-through select operator MUX_1151_inst
    position_buffer <= CONCAT_u1_u5_1144_wire when (found_upper_1135(0) /=  '0') else MUX_1150_wire;
    -- flow-through slice operator slice_1126_inst
    fp_16_upper_1127 <= fp_32_buffer(31 downto 16);
    -- flow-through slice operator slice_1130_inst
    fp_16_lower_1131 <= fp_32_buffer(15 downto 0);
    -- flow through binary operator CONCAT_u1_u5_1144_inst
    process(R_ONE_1_1142_wire_constant, fp_16_upper_index_1135) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_1142_wire_constant, fp_16_upper_index_1135, tmp_var);
      CONCAT_u1_u5_1144_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u5_1148_inst
    process(R_ZERO_1_1146_wire_constant, fp_16_lower_index_1139) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_1_1146_wire_constant, fp_16_lower_index_1139, tmp_var);
      CONCAT_u1_u5_1148_wire <= tmp_var; --
    end process;
    -- flow through binary operator OR_u1_u1_1156_inst
    found_buffer <= (found_upper_1135 or found_lower_1139);
    volatile_operator_find_left_16_799: find_left_16_Volatile port map(fp_16 => fp_16_upper_1127, position => fp_16_upper_index_1135, found => found_upper_1135); 
    volatile_operator_find_left_16_800: find_left_16_Volatile port map(fp_16 => fp_16_lower_1131, position => fp_16_lower_index_1139, found => found_lower_1139); 
    -- 
  end Block; -- data_path
  -- 
end find_left_32_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity find_left_4_Volatile is -- 
  port ( -- 
    fp_4 : in  std_logic_vector(3 downto 0);
    position : out  std_logic_vector(1 downto 0);
    found : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity find_left_4_Volatile;
architecture find_left_4_Volatile_arch of find_left_4_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(4-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal fp_4_buffer :  std_logic_vector(3 downto 0);
  -- output port buffer signals
  signal position_buffer :  std_logic_vector(1 downto 0);
  signal found_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  fp_4_buffer <= fp_4;
  -- output handling  -------------------------------------------------------
  position <= position_buffer;
  found <= found_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1033_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1032_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1017_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1020_wire : std_logic_vector(0 downto 0);
    signal x0_1013 : std_logic_vector(0 downto 0);
    signal x1_1009 : std_logic_vector(0 downto 0);
    signal x2_1005 : std_logic_vector(0 downto 0);
    signal x3_1001 : std_logic_vector(0 downto 0);
    signal y0_1035 : std_logic_vector(0 downto 0);
    signal y1_1027 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_1000_inst
    x3_1001 <= fp_4_buffer(3 downto 3);
    -- flow-through slice operator slice_1004_inst
    x2_1005 <= fp_4_buffer(2 downto 2);
    -- flow-through slice operator slice_1008_inst
    x1_1009 <= fp_4_buffer(1 downto 1);
    -- flow-through slice operator slice_1012_inst
    x0_1013 <= fp_4_buffer(0 downto 0);
    -- flow through binary operator AND_u1_u1_1033_inst
    AND_u1_u1_1033_wire <= (x1_1009 and NOT_u1_u1_1032_wire);
    -- flow through binary operator CONCAT_u1_u2_1039_inst
    process(y1_1027, y0_1035) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(y1_1027, y0_1035, tmp_var);
      position_buffer <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1032_inst
    process(x2_1005) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", x2_1005, tmp_var);
      NOT_u1_u1_1032_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_1017_inst
    OR_u1_u1_1017_wire <= (x3_1001 or x2_1005);
    -- flow through binary operator OR_u1_u1_1020_inst
    OR_u1_u1_1020_wire <= (x1_1009 or x0_1013);
    -- flow through binary operator OR_u1_u1_1021_inst
    found_buffer <= (OR_u1_u1_1017_wire or OR_u1_u1_1020_wire);
    -- flow through binary operator OR_u1_u1_1026_inst
    y1_1027 <= (x3_1001 or x2_1005);
    -- flow through binary operator OR_u1_u1_1034_inst
    y0_1035 <= (x3_1001 or AND_u1_u1_1033_wire);
    -- 
  end Block; -- data_path
  -- 
end find_left_4_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity find_left_8_Volatile is -- 
  port ( -- 
    fp_8 : in  std_logic_vector(7 downto 0);
    position : out  std_logic_vector(2 downto 0);
    found : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity find_left_8_Volatile;
architecture find_left_8_Volatile_arch of find_left_8_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal fp_8_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal position_buffer :  std_logic_vector(2 downto 0);
  signal found_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  component find_left_4_Volatile is -- 
    port ( -- 
      fp_4 : in  std_logic_vector(3 downto 0);
      position : out  std_logic_vector(1 downto 0);
      found : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  fp_8_buffer <= fp_8;
  -- output handling  -------------------------------------------------------
  position <= position_buffer;
  found <= found_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u3_1066_wire : std_logic_vector(2 downto 0);
    signal CONCAT_u1_u3_1070_wire : std_logic_vector(2 downto 0);
    signal MUX_1072_wire : std_logic_vector(2 downto 0);
    signal R_ONE_1_1064_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_1068_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_3_1071_wire_constant : std_logic_vector(2 downto 0);
    signal found_lower_1061 : std_logic_vector(0 downto 0);
    signal found_upper_1057 : std_logic_vector(0 downto 0);
    signal fp_4_lower_1053 : std_logic_vector(3 downto 0);
    signal fp_4_lower_index_1061 : std_logic_vector(1 downto 0);
    signal fp_4_upper_1049 : std_logic_vector(3 downto 0);
    signal fp_4_upper_index_1057 : std_logic_vector(1 downto 0);
    -- 
  begin -- 
    R_ONE_1_1064_wire_constant <= "1";
    R_ZERO_1_1068_wire_constant <= "0";
    R_ZERO_3_1071_wire_constant <= "000";
    -- flow-through select operator MUX_1072_inst
    MUX_1072_wire <= CONCAT_u1_u3_1070_wire when (found_lower_1061(0) /=  '0') else R_ZERO_3_1071_wire_constant;
    -- flow-through select operator MUX_1073_inst
    position_buffer <= CONCAT_u1_u3_1066_wire when (found_upper_1057(0) /=  '0') else MUX_1072_wire;
    -- flow-through slice operator slice_1048_inst
    fp_4_upper_1049 <= fp_8_buffer(7 downto 4);
    -- flow-through slice operator slice_1052_inst
    fp_4_lower_1053 <= fp_8_buffer(3 downto 0);
    -- flow through binary operator CONCAT_u1_u3_1066_inst
    process(R_ONE_1_1064_wire_constant, fp_4_upper_index_1057) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_1064_wire_constant, fp_4_upper_index_1057, tmp_var);
      CONCAT_u1_u3_1066_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u3_1070_inst
    process(R_ZERO_1_1068_wire_constant, fp_4_lower_index_1061) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_1_1068_wire_constant, fp_4_lower_index_1061, tmp_var);
      CONCAT_u1_u3_1070_wire <= tmp_var; --
    end process;
    -- flow through binary operator OR_u1_u1_1078_inst
    found_buffer <= (found_upper_1057 or found_lower_1061);
    volatile_operator_find_left_4_735: find_left_4_Volatile port map(fp_4 => fp_4_upper_1049, position => fp_4_upper_index_1057, found => found_upper_1057); 
    volatile_operator_find_left_4_736: find_left_4_Volatile port map(fp_4 => fp_4_lower_1053, position => fp_4_lower_index_1061, found => found_lower_1061); 
    -- 
  end Block; -- data_path
  -- 
end find_left_8_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity find_leftmost_64_Volatile is -- 
  port ( -- 
    fp_64 : in  std_logic_vector(63 downto 0);
    position : out  std_logic_vector(5 downto 0);
    found : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity find_leftmost_64_Volatile;
architecture find_leftmost_64_Volatile_arch of find_leftmost_64_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(64-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal fp_64_buffer :  std_logic_vector(63 downto 0);
  -- output port buffer signals
  signal position_buffer :  std_logic_vector(5 downto 0);
  signal found_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  component find_left_32_Volatile is -- 
    port ( -- 
      fp_32 : in  std_logic_vector(31 downto 0);
      position : out  std_logic_vector(4 downto 0);
      found : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  fp_64_buffer <= fp_64;
  -- output handling  -------------------------------------------------------
  position <= position_buffer;
  found <= found_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u6_1183_wire : std_logic_vector(5 downto 0);
    signal CONCAT_u1_u6_1187_wire : std_logic_vector(5 downto 0);
    signal MUX_1189_wire : std_logic_vector(5 downto 0);
    signal R_ONE_1_1181_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_1185_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_6_1188_wire_constant : std_logic_vector(5 downto 0);
    signal found_lower_1178 : std_logic_vector(0 downto 0);
    signal found_upper_1174 : std_logic_vector(0 downto 0);
    signal fp_32_lower_1170 : std_logic_vector(31 downto 0);
    signal fp_32_lower_index_1178 : std_logic_vector(4 downto 0);
    signal fp_32_upper_1166 : std_logic_vector(31 downto 0);
    signal fp_32_upper_index_1174 : std_logic_vector(4 downto 0);
    -- 
  begin -- 
    R_ONE_1_1181_wire_constant <= "1";
    R_ZERO_1_1185_wire_constant <= "0";
    R_ZERO_6_1188_wire_constant <= "000000";
    -- flow-through select operator MUX_1189_inst
    MUX_1189_wire <= CONCAT_u1_u6_1187_wire when (found_lower_1178(0) /=  '0') else R_ZERO_6_1188_wire_constant;
    -- flow-through select operator MUX_1190_inst
    position_buffer <= CONCAT_u1_u6_1183_wire when (found_upper_1174(0) /=  '0') else MUX_1189_wire;
    -- flow-through slice operator slice_1165_inst
    fp_32_upper_1166 <= fp_64_buffer(63 downto 32);
    -- flow-through slice operator slice_1169_inst
    fp_32_lower_1170 <= fp_64_buffer(31 downto 0);
    -- flow through binary operator CONCAT_u1_u6_1183_inst
    process(R_ONE_1_1181_wire_constant, fp_32_upper_index_1174) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_1181_wire_constant, fp_32_upper_index_1174, tmp_var);
      CONCAT_u1_u6_1183_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u6_1187_inst
    process(R_ZERO_1_1185_wire_constant, fp_32_lower_index_1178) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_1_1185_wire_constant, fp_32_lower_index_1178, tmp_var);
      CONCAT_u1_u6_1187_wire <= tmp_var; --
    end process;
    -- flow through binary operator OR_u1_u1_1195_inst
    found_buffer <= (found_upper_1174 or found_lower_1178);
    volatile_operator_find_left_32_831: find_left_32_Volatile port map(fp_32 => fp_32_upper_1166, position => fp_32_upper_index_1174, found => found_upper_1174); 
    volatile_operator_find_left_32_832: find_left_32_Volatile port map(fp_32 => fp_32_lower_1170, position => fp_32_lower_index_1178, found => found_lower_1178); 
    -- 
  end Block; -- data_path
  -- 
end find_leftmost_64_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity i32_add_sub_Volatile is -- 
  port ( -- 
    subtract_flag : in  std_logic_vector(0 downto 0);
    with_carry : in  std_logic_vector(0 downto 0);
    set_cc : in  std_logic_vector(0 downto 0);
    tagged_op : in  std_logic_vector(0 downto 0);
    trap_on_ovflow : in  std_logic_vector(0 downto 0);
    Ni : in  std_logic_vector(0 downto 0);
    Zi : in  std_logic_vector(0 downto 0);
    Vi : in  std_logic_vector(0 downto 0);
    Ci : in  std_logic_vector(0 downto 0);
    x : in  std_logic_vector(31 downto 0);
    y : in  std_logic_vector(31 downto 0);
    result : out  std_logic_vector(31 downto 0);
    No : out  std_logic_vector(0 downto 0);
    Zo : out  std_logic_vector(0 downto 0);
    Vo : out  std_logic_vector(0 downto 0);
    Co : out  std_logic_vector(0 downto 0);
    overflow_trap : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity i32_add_sub_Volatile;
architecture i32_add_sub_Volatile_arch of i32_add_sub_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(73-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal subtract_flag_buffer :  std_logic_vector(0 downto 0);
  signal with_carry_buffer :  std_logic_vector(0 downto 0);
  signal set_cc_buffer :  std_logic_vector(0 downto 0);
  signal tagged_op_buffer :  std_logic_vector(0 downto 0);
  signal trap_on_ovflow_buffer :  std_logic_vector(0 downto 0);
  signal Ni_buffer :  std_logic_vector(0 downto 0);
  signal Zi_buffer :  std_logic_vector(0 downto 0);
  signal Vi_buffer :  std_logic_vector(0 downto 0);
  signal Ci_buffer :  std_logic_vector(0 downto 0);
  signal x_buffer :  std_logic_vector(31 downto 0);
  signal y_buffer :  std_logic_vector(31 downto 0);
  -- output port buffer signals
  signal result_buffer :  std_logic_vector(31 downto 0);
  signal No_buffer :  std_logic_vector(0 downto 0);
  signal Zo_buffer :  std_logic_vector(0 downto 0);
  signal Vo_buffer :  std_logic_vector(0 downto 0);
  signal Co_buffer :  std_logic_vector(0 downto 0);
  signal overflow_trap_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  subtract_flag_buffer <= subtract_flag;
  with_carry_buffer <= with_carry;
  set_cc_buffer <= set_cc;
  tagged_op_buffer <= tagged_op;
  trap_on_ovflow_buffer <= trap_on_ovflow;
  Ni_buffer <= Ni;
  Zi_buffer <= Zi;
  Vi_buffer <= Vi;
  Ci_buffer <= Ci;
  x_buffer <= x;
  y_buffer <= y;
  -- output handling  -------------------------------------------------------
  result <= result_buffer;
  No <= No_buffer;
  Zo <= Zo_buffer;
  Vo <= Vo_buffer;
  Co <= Co_buffer;
  overflow_trap <= overflow_trap_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_6813_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6817_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6846_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6851_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6860_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6864_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6875_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6880_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6888_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6892_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6911_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6917_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6965_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6977_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_6991_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7003_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6842_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6845_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6849_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6854_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6858_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6863_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6870_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6873_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6878_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6883_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6887_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6891_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6936_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6961_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6964_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6968_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6972_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6975_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6986_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6990_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6994_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_6997_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_7001_wire : std_logic_vector(0 downto 0);
    signal Co_add_6981 : std_logic_vector(0 downto 0);
    signal Co_sub_7007 : std_logic_vector(0 downto 0);
    signal EQ_u32_u1_6944_wire : std_logic_vector(0 downto 0);
    signal MUX_6953_wire : std_logic_vector(0 downto 0);
    signal NEQ_u2_u1_6906_wire : std_logic_vector(0 downto 0);
    signal NEQ_u2_u1_6910_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6814_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6850_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6855_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6859_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6874_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6879_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6884_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6926_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6969_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6987_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_6998_wire : std_logic_vector(0 downto 0);
    signal NOT_u32_u32_6805_wire : std_logic_vector(31 downto 0);
    signal OR_u1_u1_6924_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6976_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_6978_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_7002_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_7004_wire : std_logic_vector(0 downto 0);
    signal add_one_6819 : std_logic_vector(0 downto 0);
    signal konst_6841_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6844_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6848_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6853_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6857_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6862_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6869_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6872_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6877_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6882_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6886_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6890_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6905_wire_constant : std_logic_vector(1 downto 0);
    signal konst_6909_wire_constant : std_logic_vector(1 downto 0);
    signal konst_6935_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6943_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6960_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6963_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6967_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6971_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6974_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6985_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6989_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6993_wire_constant : std_logic_vector(31 downto 0);
    signal konst_6996_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7000_wire_constant : std_logic_vector(31 downto 0);
    signal op_2_6808 : std_logic_vector(31 downto 0);
    signal overflow_trap_raw_6920 : std_logic_vector(0 downto 0);
    signal raw_result_6838 : std_logic_vector(31 downto 0);
    signal slice_6904_wire : std_logic_vector(1 downto 0);
    signal slice_6908_wire : std_logic_vector(1 downto 0);
    signal sum_33_6834 : std_logic_vector(32 downto 0);
    signal sum_operand_1_6824 : std_logic_vector(32 downto 0);
    signal sum_operand_2_6829 : std_logic_vector(32 downto 0);
    signal tV_6900 : std_logic_vector(0 downto 0);
    signal tV_add_6866 : std_logic_vector(0 downto 0);
    signal tV_sub_6894 : std_logic_vector(0 downto 0);
    signal tag_tV_6913 : std_logic_vector(0 downto 0);
    signal update_flags_6928 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_6841_wire_constant <= "00000000000000000000000000011111";
    konst_6844_wire_constant <= "00000000000000000000000000011111";
    konst_6848_wire_constant <= "00000000000000000000000000011111";
    konst_6853_wire_constant <= "00000000000000000000000000011111";
    konst_6857_wire_constant <= "00000000000000000000000000011111";
    konst_6862_wire_constant <= "00000000000000000000000000011111";
    konst_6869_wire_constant <= "00000000000000000000000000011111";
    konst_6872_wire_constant <= "00000000000000000000000000011111";
    konst_6877_wire_constant <= "00000000000000000000000000011111";
    konst_6882_wire_constant <= "00000000000000000000000000011111";
    konst_6886_wire_constant <= "00000000000000000000000000011111";
    konst_6890_wire_constant <= "00000000000000000000000000011111";
    konst_6905_wire_constant <= "00";
    konst_6909_wire_constant <= "00";
    konst_6935_wire_constant <= "00000000000000000000000000011111";
    konst_6943_wire_constant <= "00000000000000000000000000000000";
    konst_6960_wire_constant <= "00000000000000000000000000011111";
    konst_6963_wire_constant <= "00000000000000000000000000011111";
    konst_6967_wire_constant <= "00000000000000000000000000011111";
    konst_6971_wire_constant <= "00000000000000000000000000011111";
    konst_6974_wire_constant <= "00000000000000000000000000011111";
    konst_6985_wire_constant <= "00000000000000000000000000011111";
    konst_6989_wire_constant <= "00000000000000000000000000011111";
    konst_6993_wire_constant <= "00000000000000000000000000011111";
    konst_6996_wire_constant <= "00000000000000000000000000011111";
    konst_7000_wire_constant <= "00000000000000000000000000011111";
    -- flow-through select operator MUX_6807_inst
    op_2_6808 <= NOT_u32_u32_6805_wire when (subtract_flag_buffer(0) /=  '0') else y_buffer;
    -- flow-through select operator MUX_6818_inst
    add_one_6819 <= NOT_u1_u1_6814_wire when (subtract_flag_buffer(0) /=  '0') else AND_u1_u1_6817_wire;
    -- flow-through select operator MUX_6899_inst
    tV_6900 <= tV_sub_6894 when (subtract_flag_buffer(0) /=  '0') else tV_add_6866;
    -- flow-through select operator MUX_6938_inst
    No_buffer <= BITSEL_u32_u1_6936_wire when (update_flags_6928(0) /=  '0') else Ni_buffer;
    -- flow-through select operator MUX_6946_inst
    Zo_buffer <= EQ_u32_u1_6944_wire when (update_flags_6928(0) /=  '0') else Zi_buffer;
    -- flow-through select operator MUX_6953_inst
    MUX_6953_wire <= tag_tV_6913 when (tagged_op_buffer(0) /=  '0') else tV_6900;
    -- flow-through select operator MUX_6955_inst
    Vo_buffer <= MUX_6953_wire when (update_flags_6928(0) /=  '0') else Vi_buffer;
    -- flow-through select operator MUX_6980_inst
    Co_add_6981 <= OR_u1_u1_6978_wire when (update_flags_6928(0) /=  '0') else Ci_buffer;
    -- flow-through select operator MUX_7006_inst
    Co_sub_7007 <= OR_u1_u1_7004_wire when (update_flags_6928(0) /=  '0') else Ci_buffer;
    -- flow-through select operator MUX_7012_inst
    Co_buffer <= Co_sub_7007 when (subtract_flag_buffer(0) /=  '0') else Co_add_6981;
    -- flow-through slice operator slice_6837_inst
    raw_result_6838 <= sum_33_6834(32 downto 1);
    -- flow-through slice operator slice_6904_inst
    slice_6904_wire <= x_buffer(1 downto 0);
    -- flow-through slice operator slice_6908_inst
    slice_6908_wire <= y_buffer(1 downto 0);
    -- interlock W_overflow_trap_6929_inst
    process(overflow_trap_raw_6920) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := overflow_trap_raw_6920(0 downto 0);
      overflow_trap_buffer <= tmp_var; -- 
    end process;
    -- interlock W_result_7014_inst
    process(raw_result_6838) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := raw_result_6838(31 downto 0);
      result_buffer <= tmp_var; -- 
    end process;
    -- flow through binary operator ADD_u33_u33_6833_inst
    sum_33_6834 <= std_logic_vector(unsigned(sum_operand_1_6824) + unsigned(sum_operand_2_6829));
    -- flow through binary operator AND_u1_u1_6813_inst
    AND_u1_u1_6813_wire <= (Ci_buffer and with_carry_buffer);
    -- flow through binary operator AND_u1_u1_6817_inst
    AND_u1_u1_6817_wire <= (Ci_buffer and with_carry_buffer);
    -- flow through binary operator AND_u1_u1_6846_inst
    AND_u1_u1_6846_wire <= (BITSEL_u32_u1_6842_wire and BITSEL_u32_u1_6845_wire);
    -- flow through binary operator AND_u1_u1_6851_inst
    AND_u1_u1_6851_wire <= (AND_u1_u1_6846_wire and NOT_u1_u1_6850_wire);
    -- flow through binary operator AND_u1_u1_6860_inst
    AND_u1_u1_6860_wire <= (NOT_u1_u1_6855_wire and NOT_u1_u1_6859_wire);
    -- flow through binary operator AND_u1_u1_6864_inst
    AND_u1_u1_6864_wire <= (AND_u1_u1_6860_wire and BITSEL_u32_u1_6863_wire);
    -- flow through binary operator AND_u1_u1_6875_inst
    AND_u1_u1_6875_wire <= (BITSEL_u32_u1_6870_wire and NOT_u1_u1_6874_wire);
    -- flow through binary operator AND_u1_u1_6880_inst
    AND_u1_u1_6880_wire <= (AND_u1_u1_6875_wire and NOT_u1_u1_6879_wire);
    -- flow through binary operator AND_u1_u1_6888_inst
    AND_u1_u1_6888_wire <= (NOT_u1_u1_6884_wire and BITSEL_u32_u1_6887_wire);
    -- flow through binary operator AND_u1_u1_6892_inst
    AND_u1_u1_6892_wire <= (AND_u1_u1_6888_wire and BITSEL_u32_u1_6891_wire);
    -- flow through binary operator AND_u1_u1_6911_inst
    AND_u1_u1_6911_wire <= (NEQ_u2_u1_6906_wire and NEQ_u2_u1_6910_wire);
    -- flow through binary operator AND_u1_u1_6917_inst
    AND_u1_u1_6917_wire <= (tagged_op_buffer and tag_tV_6913);
    -- flow through binary operator AND_u1_u1_6919_inst
    overflow_trap_raw_6920 <= (AND_u1_u1_6917_wire and trap_on_ovflow_buffer);
    -- flow through binary operator AND_u1_u1_6927_inst
    update_flags_6928 <= (OR_u1_u1_6924_wire and NOT_u1_u1_6926_wire);
    -- flow through binary operator AND_u1_u1_6965_inst
    AND_u1_u1_6965_wire <= (BITSEL_u32_u1_6961_wire and BITSEL_u32_u1_6964_wire);
    -- flow through binary operator AND_u1_u1_6977_inst
    AND_u1_u1_6977_wire <= (NOT_u1_u1_6969_wire and OR_u1_u1_6976_wire);
    -- flow through binary operator AND_u1_u1_6991_inst
    AND_u1_u1_6991_wire <= (NOT_u1_u1_6987_wire and BITSEL_u32_u1_6990_wire);
    -- flow through binary operator AND_u1_u1_7003_inst
    AND_u1_u1_7003_wire <= (BITSEL_u32_u1_6994_wire and OR_u1_u1_7002_wire);
    -- flow through binary operator BITSEL_u32_u1_6842_inst
    process(x_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(x_buffer, konst_6841_wire_constant, tmp_var);
      BITSEL_u32_u1_6842_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6845_inst
    process(y_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(y_buffer, konst_6844_wire_constant, tmp_var);
      BITSEL_u32_u1_6845_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6849_inst
    process(raw_result_6838) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(raw_result_6838, konst_6848_wire_constant, tmp_var);
      BITSEL_u32_u1_6849_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6854_inst
    process(x_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(x_buffer, konst_6853_wire_constant, tmp_var);
      BITSEL_u32_u1_6854_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6858_inst
    process(y_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(y_buffer, konst_6857_wire_constant, tmp_var);
      BITSEL_u32_u1_6858_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6863_inst
    process(raw_result_6838) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(raw_result_6838, konst_6862_wire_constant, tmp_var);
      BITSEL_u32_u1_6863_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6870_inst
    process(x_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(x_buffer, konst_6869_wire_constant, tmp_var);
      BITSEL_u32_u1_6870_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6873_inst
    process(y_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(y_buffer, konst_6872_wire_constant, tmp_var);
      BITSEL_u32_u1_6873_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6878_inst
    process(raw_result_6838) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(raw_result_6838, konst_6877_wire_constant, tmp_var);
      BITSEL_u32_u1_6878_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6883_inst
    process(x_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(x_buffer, konst_6882_wire_constant, tmp_var);
      BITSEL_u32_u1_6883_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6887_inst
    process(y_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(y_buffer, konst_6886_wire_constant, tmp_var);
      BITSEL_u32_u1_6887_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6891_inst
    process(raw_result_6838) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(raw_result_6838, konst_6890_wire_constant, tmp_var);
      BITSEL_u32_u1_6891_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6936_inst
    process(raw_result_6838) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(raw_result_6838, konst_6935_wire_constant, tmp_var);
      BITSEL_u32_u1_6936_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6961_inst
    process(x_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(x_buffer, konst_6960_wire_constant, tmp_var);
      BITSEL_u32_u1_6961_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6964_inst
    process(y_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(y_buffer, konst_6963_wire_constant, tmp_var);
      BITSEL_u32_u1_6964_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6968_inst
    process(raw_result_6838) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(raw_result_6838, konst_6967_wire_constant, tmp_var);
      BITSEL_u32_u1_6968_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6972_inst
    process(x_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(x_buffer, konst_6971_wire_constant, tmp_var);
      BITSEL_u32_u1_6972_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6975_inst
    process(y_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(y_buffer, konst_6974_wire_constant, tmp_var);
      BITSEL_u32_u1_6975_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6986_inst
    process(x_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(x_buffer, konst_6985_wire_constant, tmp_var);
      BITSEL_u32_u1_6986_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6990_inst
    process(y_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(y_buffer, konst_6989_wire_constant, tmp_var);
      BITSEL_u32_u1_6990_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6994_inst
    process(raw_result_6838) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(raw_result_6838, konst_6993_wire_constant, tmp_var);
      BITSEL_u32_u1_6994_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_6997_inst
    process(x_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(x_buffer, konst_6996_wire_constant, tmp_var);
      BITSEL_u32_u1_6997_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_7001_inst
    process(y_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(y_buffer, konst_7000_wire_constant, tmp_var);
      BITSEL_u32_u1_7001_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u32_u33_6823_inst
    process(x_buffer, add_one_6819) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(x_buffer, add_one_6819, tmp_var);
      sum_operand_1_6824 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u32_u33_6828_inst
    process(op_2_6808, add_one_6819) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(op_2_6808, add_one_6819, tmp_var);
      sum_operand_2_6829 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_6944_inst
    process(raw_result_6838) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(raw_result_6838, konst_6943_wire_constant, tmp_var);
      EQ_u32_u1_6944_wire <= tmp_var; --
    end process;
    -- flow through binary operator NEQ_u2_u1_6906_inst
    process(slice_6904_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(slice_6904_wire, konst_6905_wire_constant, tmp_var);
      NEQ_u2_u1_6906_wire <= tmp_var; --
    end process;
    -- flow through binary operator NEQ_u2_u1_6910_inst
    process(slice_6908_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(slice_6908_wire, konst_6909_wire_constant, tmp_var);
      NEQ_u2_u1_6910_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_6814_inst
    process(AND_u1_u1_6813_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", AND_u1_u1_6813_wire, tmp_var);
      NOT_u1_u1_6814_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6850_inst
    process(BITSEL_u32_u1_6849_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_6849_wire, tmp_var);
      NOT_u1_u1_6850_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6855_inst
    process(BITSEL_u32_u1_6854_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_6854_wire, tmp_var);
      NOT_u1_u1_6855_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6859_inst
    process(BITSEL_u32_u1_6858_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_6858_wire, tmp_var);
      NOT_u1_u1_6859_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6874_inst
    process(BITSEL_u32_u1_6873_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_6873_wire, tmp_var);
      NOT_u1_u1_6874_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6879_inst
    process(BITSEL_u32_u1_6878_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_6878_wire, tmp_var);
      NOT_u1_u1_6879_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6884_inst
    process(BITSEL_u32_u1_6883_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_6883_wire, tmp_var);
      NOT_u1_u1_6884_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6926_inst
    process(overflow_trap_raw_6920) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", overflow_trap_raw_6920, tmp_var);
      NOT_u1_u1_6926_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6969_inst
    process(BITSEL_u32_u1_6968_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_6968_wire, tmp_var);
      NOT_u1_u1_6969_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6987_inst
    process(BITSEL_u32_u1_6986_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_6986_wire, tmp_var);
      NOT_u1_u1_6987_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_6998_inst
    process(BITSEL_u32_u1_6997_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_6997_wire, tmp_var);
      NOT_u1_u1_6998_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u32_u32_6805_inst
    process(y_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", y_buffer, tmp_var);
      NOT_u32_u32_6805_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_6865_inst
    tV_add_6866 <= (AND_u1_u1_6851_wire or AND_u1_u1_6864_wire);
    -- flow through binary operator OR_u1_u1_6893_inst
    tV_sub_6894 <= (AND_u1_u1_6880_wire or AND_u1_u1_6892_wire);
    -- flow through binary operator OR_u1_u1_6912_inst
    tag_tV_6913 <= (tV_6900 or AND_u1_u1_6911_wire);
    -- flow through binary operator OR_u1_u1_6924_inst
    OR_u1_u1_6924_wire <= (tagged_op_buffer or set_cc_buffer);
    -- flow through binary operator OR_u1_u1_6976_inst
    OR_u1_u1_6976_wire <= (BITSEL_u32_u1_6972_wire or BITSEL_u32_u1_6975_wire);
    -- flow through binary operator OR_u1_u1_6978_inst
    OR_u1_u1_6978_wire <= (AND_u1_u1_6965_wire or AND_u1_u1_6977_wire);
    -- flow through binary operator OR_u1_u1_7002_inst
    OR_u1_u1_7002_wire <= (NOT_u1_u1_6998_wire or BITSEL_u32_u1_7001_wire);
    -- flow through binary operator OR_u1_u1_7004_inst
    OR_u1_u1_7004_wire <= (AND_u1_u1_6991_wire or AND_u1_u1_7003_wire);
    -- 
  end Block; -- data_path
  -- 
end i32_add_sub_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity i32_div is -- 
  generic (tag_length : integer); 
  port ( -- 
    signed_div : in  std_logic_vector(0 downto 0);
    set_cc : in  std_logic_vector(0 downto 0);
    y_in : in  std_logic_vector(31 downto 0);
    dividend : in  std_logic_vector(31 downto 0);
    divisor : in  std_logic_vector(31 downto 0);
    result : out  std_logic_vector(31 downto 0);
    No : out  std_logic_vector(0 downto 0);
    Zo : out  std_logic_vector(0 downto 0);
    Vo : out  std_logic_vector(0 downto 0);
    Co : out  std_logic_vector(0 downto 0);
    u64_true_divide_revised_call_reqs : out  std_logic_vector(0 downto 0);
    u64_true_divide_revised_call_acks : in   std_logic_vector(0 downto 0);
    u64_true_divide_revised_call_data : out  std_logic_vector(95 downto 0);
    u64_true_divide_revised_call_tag  :  out  std_logic_vector(0 downto 0);
    u64_true_divide_revised_return_reqs : out  std_logic_vector(0 downto 0);
    u64_true_divide_revised_return_acks : in   std_logic_vector(0 downto 0);
    u64_true_divide_revised_return_data : in   std_logic_vector(63 downto 0);
    u64_true_divide_revised_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity i32_div;
architecture i32_div_arch of i32_div is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 98)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal signed_div_buffer :  std_logic_vector(0 downto 0);
  signal signed_div_update_enable: Boolean;
  signal set_cc_buffer :  std_logic_vector(0 downto 0);
  signal set_cc_update_enable: Boolean;
  signal y_in_buffer :  std_logic_vector(31 downto 0);
  signal y_in_update_enable: Boolean;
  signal dividend_buffer :  std_logic_vector(31 downto 0);
  signal dividend_update_enable: Boolean;
  signal divisor_buffer :  std_logic_vector(31 downto 0);
  signal divisor_update_enable: Boolean;
  -- output port buffer signals
  signal result_buffer :  std_logic_vector(31 downto 0);
  signal result_update_enable: Boolean;
  signal No_buffer :  std_logic_vector(0 downto 0);
  signal No_update_enable: Boolean;
  signal Zo_buffer :  std_logic_vector(0 downto 0);
  signal Zo_update_enable: Boolean;
  signal Vo_buffer :  std_logic_vector(0 downto 0);
  signal Vo_update_enable: Boolean;
  signal Co_buffer :  std_logic_vector(0 downto 0);
  signal i32_div_CP_774_start: Boolean;
  signal i32_div_CP_774_symbol: Boolean;
  -- volatile/operator module components. 
  component u_cmp_32_Volatile is -- 
    port ( -- 
      a : in  std_logic_vector(31 downto 0);
      b : in  std_logic_vector(31 downto 0);
      l : out  std_logic_vector(0 downto 0);
      g : out  std_logic_vector(0 downto 0);
      e : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component twos_complement_64_Volatile is -- 
    port ( -- 
      A : in  std_logic_vector(63 downto 0);
      B : out  std_logic_vector(63 downto 0)-- 
    );
    -- 
  end component; 
  component u64_true_divide_revised is -- 
    generic (tag_length : integer); 
    port ( -- 
      udividend : in  std_logic_vector(63 downto 0);
      udivisor : in  std_logic_vector(31 downto 0);
      quotient : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component twos_complement_32_Volatile is -- 
    port ( -- 
      A : in  std_logic_vector(31 downto 0);
      B : out  std_logic_vector(31 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal W_Vo_7777_inst_req_0 : boolean;
  signal EQ_u32_u1_7775_inst_ack_0 : boolean;
  signal EQ_u32_u1_7775_inst_req_0 : boolean;
  signal W_Vo_7777_inst_ack_1 : boolean;
  signal W_Vo_7777_inst_req_1 : boolean;
  signal EQ_u32_u1_7775_inst_req_1 : boolean;
  signal W_Vo_7777_inst_ack_0 : boolean;
  signal EQ_u32_u1_7775_inst_ack_1 : boolean;
  signal BITSEL_u32_u1_7770_inst_ack_1 : boolean;
  signal BITSEL_u32_u1_7770_inst_req_1 : boolean;
  signal BITSEL_u32_u1_7770_inst_ack_0 : boolean;
  signal BITSEL_u32_u1_7770_inst_req_0 : boolean;
  signal W_result_7764_inst_ack_1 : boolean;
  signal W_result_7764_inst_req_1 : boolean;
  signal W_result_7764_inst_ack_0 : boolean;
  signal W_result_7764_inst_req_0 : boolean;
  signal call_stmt_7685_call_ack_1 : boolean;
  signal call_stmt_7685_call_req_1 : boolean;
  signal call_stmt_7685_call_ack_0 : boolean;
  signal call_stmt_7685_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "i32_div_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 98) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= signed_div;
  signed_div_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(1 downto 1) <= set_cc;
  set_cc_buffer <= in_buffer_data_out(1 downto 1);
  in_buffer_data_in(33 downto 2) <= y_in;
  y_in_buffer <= in_buffer_data_out(33 downto 2);
  in_buffer_data_in(65 downto 34) <= dividend;
  dividend_buffer <= in_buffer_data_out(65 downto 34);
  in_buffer_data_in(97 downto 66) <= divisor;
  divisor_buffer <= in_buffer_data_out(97 downto 66);
  in_buffer_data_in(tag_length + 97 downto 98) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 97 downto 98);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  i32_div_CP_774_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "i32_div_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 36) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= result_buffer;
  result <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(32 downto 32) <= No_buffer;
  No <= out_buffer_data_out(32 downto 32);
  out_buffer_data_in(33 downto 33) <= Zo_buffer;
  Zo <= out_buffer_data_out(33 downto 33);
  out_buffer_data_in(34 downto 34) <= Vo_buffer;
  Vo <= out_buffer_data_out(34 downto 34);
  Co_buffer <= "0";
  out_buffer_data_in(35 downto 35) <= Co_buffer;
  Co <= out_buffer_data_out(35 downto 35);
  out_buffer_data_in(tag_length + 35 downto 36) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 35 downto 36);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= i32_div_CP_774_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= i32_div_CP_774_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= i32_div_CP_774_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  i32_div_CP_774: Block -- control-path 
    signal i32_div_CP_774_elements: BooleanArray(11 downto 0);
    -- 
  begin -- 
    i32_div_CP_774_elements(0) <= i32_div_CP_774_start;
    i32_div_CP_774_symbol <= i32_div_CP_774_elements(11);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (20) 
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/EQ_u32_u1_7775_update_start_
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/EQ_u32_u1_7775_Update/$entry
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7779_Update/req
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/EQ_u32_u1_7775_Update/cr
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7779_update_start_
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/BITSEL_u32_u1_7770_Update/cr
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/BITSEL_u32_u1_7770_Update/$entry
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/BITSEL_u32_u1_7770_update_start_
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7779_Update/$entry
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7766_Update/req
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7766_Update/$entry
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7766_update_start_
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/call_stmt_7685_Update/ccr
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/call_stmt_7685_Update/$entry
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/call_stmt_7685_Sample/crr
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/call_stmt_7685_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/call_stmt_7685_update_start_
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/call_stmt_7685_sample_start_
      -- CP-element group 0: 	 assign_stmt_7595_to_assign_stmt_7782/$entry
      -- CP-element group 0: 	 $entry
      -- 
    req_806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => i32_div_CP_774_elements(0), ack => W_result_7764_inst_req_1); -- 
    cr_820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => i32_div_CP_774_elements(0), ack => BITSEL_u32_u1_7770_inst_req_1); -- 
    ccr_792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => i32_div_CP_774_elements(0), ack => call_stmt_7685_call_req_1); -- 
    req_848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => i32_div_CP_774_elements(0), ack => W_Vo_7777_inst_req_1); -- 
    crr_787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => i32_div_CP_774_elements(0), ack => call_stmt_7685_call_req_0); -- 
    cr_834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => i32_div_CP_774_elements(0), ack => EQ_u32_u1_7775_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_7595_to_assign_stmt_7782/call_stmt_7685_Sample/cra
      -- CP-element group 1: 	 assign_stmt_7595_to_assign_stmt_7782/call_stmt_7685_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_7595_to_assign_stmt_7782/call_stmt_7685_sample_completed_
      -- 
    cra_788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_7685_call_ack_0, ack => i32_div_CP_774_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (15) 
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7779_Sample/req
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7779_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/EQ_u32_u1_7775_Sample/rr
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/EQ_u32_u1_7775_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/EQ_u32_u1_7775_sample_start_
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/BITSEL_u32_u1_7770_Sample/rr
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/BITSEL_u32_u1_7770_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7779_sample_start_
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/BITSEL_u32_u1_7770_sample_start_
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7766_Sample/req
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7766_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7766_sample_start_
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/call_stmt_7685_Update/cca
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/call_stmt_7685_Update/$exit
      -- CP-element group 2: 	 assign_stmt_7595_to_assign_stmt_7782/call_stmt_7685_update_completed_
      -- 
    cca_793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_7685_call_ack_1, ack => i32_div_CP_774_elements(2)); -- 
    rr_815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => i32_div_CP_774_elements(2), ack => BITSEL_u32_u1_7770_inst_req_0); -- 
    req_843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => i32_div_CP_774_elements(2), ack => W_Vo_7777_inst_req_0); -- 
    req_801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => i32_div_CP_774_elements(2), ack => W_result_7764_inst_req_0); -- 
    rr_829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => i32_div_CP_774_elements(2), ack => EQ_u32_u1_7775_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7766_Sample/ack
      -- CP-element group 3: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7766_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7766_sample_completed_
      -- 
    ack_802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_result_7764_inst_ack_0, ack => i32_div_CP_774_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	11 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7766_Update/ack
      -- CP-element group 4: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7766_Update/$exit
      -- CP-element group 4: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7766_update_completed_
      -- 
    ack_807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_result_7764_inst_ack_1, ack => i32_div_CP_774_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_7595_to_assign_stmt_7782/BITSEL_u32_u1_7770_Sample/ra
      -- CP-element group 5: 	 assign_stmt_7595_to_assign_stmt_7782/BITSEL_u32_u1_7770_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_7595_to_assign_stmt_7782/BITSEL_u32_u1_7770_sample_completed_
      -- 
    ra_816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u32_u1_7770_inst_ack_0, ack => i32_div_CP_774_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	11 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_7595_to_assign_stmt_7782/BITSEL_u32_u1_7770_Update/ca
      -- CP-element group 6: 	 assign_stmt_7595_to_assign_stmt_7782/BITSEL_u32_u1_7770_Update/$exit
      -- CP-element group 6: 	 assign_stmt_7595_to_assign_stmt_7782/BITSEL_u32_u1_7770_update_completed_
      -- 
    ca_821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u32_u1_7770_inst_ack_1, ack => i32_div_CP_774_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_7595_to_assign_stmt_7782/EQ_u32_u1_7775_sample_completed_
      -- CP-element group 7: 	 assign_stmt_7595_to_assign_stmt_7782/EQ_u32_u1_7775_Sample/ra
      -- CP-element group 7: 	 assign_stmt_7595_to_assign_stmt_7782/EQ_u32_u1_7775_Sample/$exit
      -- 
    ra_830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_7775_inst_ack_0, ack => i32_div_CP_774_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	11 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_7595_to_assign_stmt_7782/EQ_u32_u1_7775_Update/$exit
      -- CP-element group 8: 	 assign_stmt_7595_to_assign_stmt_7782/EQ_u32_u1_7775_update_completed_
      -- CP-element group 8: 	 assign_stmt_7595_to_assign_stmt_7782/EQ_u32_u1_7775_Update/ca
      -- 
    ca_835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_7775_inst_ack_1, ack => i32_div_CP_774_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7779_Sample/$exit
      -- CP-element group 9: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7779_Sample/ack
      -- CP-element group 9: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7779_sample_completed_
      -- 
    ack_844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_Vo_7777_inst_ack_0, ack => i32_div_CP_774_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7779_update_completed_
      -- CP-element group 10: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7779_Update/ack
      -- CP-element group 10: 	 assign_stmt_7595_to_assign_stmt_7782/assign_stmt_7779_Update/$exit
      -- 
    ack_849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_Vo_7777_inst_ack_1, ack => i32_div_CP_774_elements(10)); -- 
    -- CP-element group 11:  join  transition  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: 	4 
    -- CP-element group 11: 	10 
    -- CP-element group 11: 	6 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 assign_stmt_7595_to_assign_stmt_7782/$exit
      -- CP-element group 11: 	 $exit
      -- 
    i32_div_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 27) := "i32_div_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= i32_div_CP_774_elements(8) & i32_div_CP_774_elements(4) & i32_div_CP_774_elements(10) & i32_div_CP_774_elements(6);
      gj_i32_div_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => i32_div_CP_774_elements(11), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_7629_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7676_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u64_u1_7749_wire : std_logic_vector(0 downto 0);
    signal EQ_u32_u1_7651_wire : std_logic_vector(0 downto 0);
    signal EQ_u32_u1_7668_wire : std_logic_vector(0 downto 0);
    signal EQ_u32_u1_7740_wire : std_logic_vector(0 downto 0);
    signal EQ_u33_u1_7730_wire : std_logic_vector(0 downto 0);
    signal EQ_u33_u1_7735_wire : std_logic_vector(0 downto 0);
    signal MUX_7619_wire : std_logic_vector(63 downto 0);
    signal MUX_7690_wire : std_logic_vector(63 downto 0);
    signal MUX_7696_wire : std_logic_vector(63 downto 0);
    signal MUX_7701_wire : std_logic_vector(63 downto 0);
    signal MUX_7722_wire : std_logic_vector(63 downto 0);
    signal MUX_7741_wire : std_logic_vector(0 downto 0);
    signal MUX_7752_wire : std_logic_vector(31 downto 0);
    signal MUX_7754_wire : std_logic_vector(31 downto 0);
    signal NOT_u1_u1_7665_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_7673_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_7675_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_7678_wire : std_logic_vector(0 downto 0);
    signal NOT_u33_u33_7734_wire_constant : std_logic_vector(32 downto 0);
    signal OR_u1_u1_7693_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_7717_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_7736_wire : std_logic_vector(0 downto 0);
    signal OR_u64_u64_7697_wire : std_logic_vector(63 downto 0);
    signal QUOTIENT_7685 : std_logic_vector(63 downto 0);
    signal R_ZERO_64_7694_wire_constant : std_logic_vector(63 downto 0);
    signal R_ZERO_64_7718_wire_constant : std_logic_vector(63 downto 0);
    signal XOR_u1_u1_7708_wire : std_logic_vector(0 downto 0);
    signal div_by_0_trap_7595 : std_logic_vector(0 downto 0);
    signal dividend_64_7605 : std_logic_vector(63 downto 0);
    signal e_7647 : std_logic_vector(0 downto 0);
    signal fQ_7724 : std_logic_vector(63 downto 0);
    signal g_7647 : std_logic_vector(0 downto 0);
    signal invert_bit_7710 : std_logic_vector(0 downto 0);
    signal inverted_dividend_64_7613 : std_logic_vector(63 downto 0);
    signal inverted_divisor_7625 : std_logic_vector(31 downto 0);
    signal inverted_no_trap_result_7713 : std_logic_vector(63 downto 0);
    signal konst_7593_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7598_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7608_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7650_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7667_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7689_wire_constant : std_logic_vector(63 downto 0);
    signal konst_7695_wire_constant : std_logic_vector(63 downto 0);
    signal konst_7700_wire_constant : std_logic_vector(63 downto 0);
    signal konst_7729_wire_constant : std_logic_vector(32 downto 0);
    signal konst_7739_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7748_wire_constant : std_logic_vector(63 downto 0);
    signal konst_7750_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7751_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7753_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7769_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7774_wire_constant : std_logic_vector(31 downto 0);
    signal l_7647 : std_logic_vector(0 downto 0);
    signal no_trap_result_7703 : std_logic_vector(63 downto 0);
    signal q_is_d_7670 : std_logic_vector(0 downto 0);
    signal run_true_divide_7680 : std_logic_vector(0 downto 0);
    signal sdividend_7600 : std_logic_vector(0 downto 0);
    signal sdivisor_7610 : std_logic_vector(0 downto 0);
    signal slice_7728_wire : std_logic_vector(32 downto 0);
    signal slice_7732_wire : std_logic_vector(32 downto 0);
    signal slice_7738_wire : std_logic_vector(31 downto 0);
    signal slice_7756_wire : std_logic_vector(31 downto 0);
    signal temp_V_7743 : std_logic_vector(0 downto 0);
    signal udividend_7622 : std_logic_vector(63 downto 0);
    signal udividend_h_7637 : std_logic_vector(31 downto 0);
    signal udividend_l_7641 : std_logic_vector(31 downto 0);
    signal udivisor_7633 : std_logic_vector(31 downto 0);
    signal vresult_7758 : std_logic_vector(31 downto 0);
    signal zero_result_7654 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u33_u33_7734_wire_constant <= "111111111111111111111111111111111";
    R_ZERO_64_7694_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    R_ZERO_64_7718_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_7593_wire_constant <= "00000000000000000000000000000000";
    konst_7598_wire_constant <= "00000000000000000000000000011111";
    konst_7608_wire_constant <= "00000000000000000000000000011111";
    konst_7650_wire_constant <= "00000000000000000000000000000000";
    konst_7667_wire_constant <= "00000000000000000000000000000001";
    konst_7689_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_7695_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_7700_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_7729_wire_constant <= "000000000000000000000000000000000";
    konst_7739_wire_constant <= "00000000000000000000000000000000";
    konst_7748_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111111";
    konst_7750_wire_constant <= "10000000000000000000000000000000";
    konst_7751_wire_constant <= "01111111111111111111111111111111";
    konst_7753_wire_constant <= "11111111111111111111111111111111";
    konst_7769_wire_constant <= "00000000000000000000000000011111";
    konst_7774_wire_constant <= "00000000000000000000000000000000";
    -- flow-through select operator MUX_7619_inst
    MUX_7619_wire <= inverted_dividend_64_7613 when (sdividend_7600(0) /=  '0') else dividend_64_7605;
    -- flow-through select operator MUX_7621_inst
    udividend_7622 <= MUX_7619_wire when (signed_div_buffer(0) /=  '0') else dividend_64_7605;
    -- flow-through select operator MUX_7632_inst
    udivisor_7633 <= inverted_divisor_7625 when (AND_u1_u1_7629_wire(0) /=  '0') else divisor_buffer;
    -- flow-through select operator MUX_7690_inst
    MUX_7690_wire <= QUOTIENT_7685 when (run_true_divide_7680(0) /=  '0') else konst_7689_wire_constant;
    -- flow-through select operator MUX_7696_inst
    MUX_7696_wire <= R_ZERO_64_7694_wire_constant when (OR_u1_u1_7693_wire(0) /=  '0') else konst_7695_wire_constant;
    -- flow-through select operator MUX_7701_inst
    MUX_7701_wire <= udividend_7622 when (q_is_d_7670(0) /=  '0') else konst_7700_wire_constant;
    -- flow-through select operator MUX_7722_inst
    MUX_7722_wire <= inverted_no_trap_result_7713 when (invert_bit_7710(0) /=  '0') else no_trap_result_7703;
    -- flow-through select operator MUX_7723_inst
    fQ_7724 <= R_ZERO_64_7718_wire_constant when (OR_u1_u1_7717_wire(0) /=  '0') else MUX_7722_wire;
    -- flow-through select operator MUX_7741_inst
    MUX_7741_wire <= OR_u1_u1_7736_wire when (signed_div_buffer(0) /=  '0') else EQ_u32_u1_7740_wire;
    -- flow-through select operator MUX_7752_inst
    MUX_7752_wire <= konst_7750_wire_constant when (BITSEL_u64_u1_7749_wire(0) /=  '0') else konst_7751_wire_constant;
    -- flow-through select operator MUX_7754_inst
    MUX_7754_wire <= MUX_7752_wire when (signed_div_buffer(0) /=  '0') else konst_7753_wire_constant;
    -- flow-through select operator MUX_7757_inst
    vresult_7758 <= MUX_7754_wire when (temp_V_7743(0) /=  '0') else slice_7756_wire;
    -- flow-through slice operator slice_7636_inst
    udividend_h_7637 <= udividend_7622(63 downto 32);
    -- flow-through slice operator slice_7640_inst
    udividend_l_7641 <= udividend_7622(31 downto 0);
    -- flow-through slice operator slice_7728_inst
    slice_7728_wire <= fQ_7724(63 downto 31);
    -- flow-through slice operator slice_7732_inst
    slice_7732_wire <= fQ_7724(63 downto 31);
    -- flow-through slice operator slice_7738_inst
    slice_7738_wire <= fQ_7724(63 downto 32);
    -- flow-through slice operator slice_7756_inst
    slice_7756_wire <= fQ_7724(31 downto 0);
    W_Vo_7777_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_Vo_7777_inst_req_0;
      W_Vo_7777_inst_ack_0<= wack(0);
      rreq(0) <= W_Vo_7777_inst_req_1;
      W_Vo_7777_inst_ack_1<= rack(0);
      W_Vo_7777_inst : InterlockBuffer generic map ( -- 
        name => "W_Vo_7777_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => temp_V_7743,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => Vo_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_result_7764_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_result_7764_inst_req_0;
      W_result_7764_inst_ack_0<= wack(0);
      rreq(0) <= W_result_7764_inst_req_1;
      W_result_7764_inst_ack_1<= rack(0);
      W_result_7764_inst : InterlockBuffer generic map ( -- 
        name => "W_result_7764_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => vresult_7758,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => result_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- flow through binary operator AND_u1_u1_7629_inst
    AND_u1_u1_7629_wire <= (signed_div_buffer and sdivisor_7610);
    -- flow through binary operator AND_u1_u1_7653_inst
    zero_result_7654 <= (EQ_u32_u1_7651_wire and l_7647);
    -- flow through binary operator AND_u1_u1_7669_inst
    q_is_d_7670 <= (NOT_u1_u1_7665_wire and EQ_u32_u1_7668_wire);
    -- flow through binary operator AND_u1_u1_7676_inst
    AND_u1_u1_7676_wire <= (NOT_u1_u1_7673_wire and NOT_u1_u1_7675_wire);
    -- flow through binary operator AND_u1_u1_7679_inst
    run_true_divide_7680 <= (AND_u1_u1_7676_wire and NOT_u1_u1_7678_wire);
    -- flow through binary operator AND_u1_u1_7709_inst
    invert_bit_7710 <= (signed_div_buffer and XOR_u1_u1_7708_wire);
    -- flow through binary operator BITSEL_u32_u1_7599_inst
    process(y_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(y_in_buffer, konst_7598_wire_constant, tmp_var);
      sdividend_7600 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_7609_inst
    process(divisor_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(divisor_buffer, konst_7608_wire_constant, tmp_var);
      sdivisor_7610 <= tmp_var; --
    end process;
    -- shared split operator group (8) : BITSEL_u32_u1_7770_inst 
    ApBitsel_group_8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= vresult_7758;
      No_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= BITSEL_u32_u1_7770_inst_req_0;
      BITSEL_u32_u1_7770_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= BITSEL_u32_u1_7770_inst_req_1;
      BITSEL_u32_u1_7770_inst_ack_1 <= ackR_unguarded(0);
      ApBitsel_group_8_gI: SplitGuardInterface generic map(name => "ApBitsel_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApBitsel",
          name => "ApBitsel_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000011111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- flow through binary operator BITSEL_u64_u1_7749_inst
    process(fQ_7724) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(fQ_7724, konst_7748_wire_constant, tmp_var);
      BITSEL_u64_u1_7749_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u32_u64_7604_inst
    process(y_in_buffer, dividend_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(y_in_buffer, dividend_buffer, tmp_var);
      dividend_64_7605 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_7594_inst
    process(divisor_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(divisor_buffer, konst_7593_wire_constant, tmp_var);
      div_by_0_trap_7595 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_7651_inst
    process(udividend_h_7637) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(udividend_h_7637, konst_7650_wire_constant, tmp_var);
      EQ_u32_u1_7651_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_7668_inst
    process(udivisor_7633) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(udivisor_7633, konst_7667_wire_constant, tmp_var);
      EQ_u32_u1_7668_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_7740_inst
    process(slice_7738_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(slice_7738_wire, konst_7739_wire_constant, tmp_var);
      EQ_u32_u1_7740_wire <= tmp_var; --
    end process;
    -- shared split operator group (15) : EQ_u32_u1_7775_inst 
    ApIntEq_group_15: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= vresult_7758;
      Zo_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u32_u1_7775_inst_req_0;
      EQ_u32_u1_7775_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_7775_inst_req_1;
      EQ_u32_u1_7775_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_15_gI: SplitGuardInterface generic map(name => "ApIntEq_group_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- flow through binary operator EQ_u33_u1_7730_inst
    process(slice_7728_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(slice_7728_wire, konst_7729_wire_constant, tmp_var);
      EQ_u33_u1_7730_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u33_u1_7735_inst
    process(slice_7732_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(slice_7732_wire, NOT_u33_u33_7734_wire_constant, tmp_var);
      EQ_u33_u1_7735_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_7665_inst
    process(zero_result_7654) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", zero_result_7654, tmp_var);
      NOT_u1_u1_7665_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_7673_inst
    process(div_by_0_trap_7595) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", div_by_0_trap_7595, tmp_var);
      NOT_u1_u1_7673_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_7675_inst
    process(zero_result_7654) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", zero_result_7654, tmp_var);
      NOT_u1_u1_7675_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_7678_inst
    process(q_is_d_7670) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", q_is_d_7670, tmp_var);
      NOT_u1_u1_7678_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_7742_inst
    process(MUX_7741_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", MUX_7741_wire, tmp_var);
      temp_V_7743 <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_7693_inst
    OR_u1_u1_7693_wire <= (div_by_0_trap_7595 or zero_result_7654);
    -- flow through binary operator OR_u1_u1_7717_inst
    OR_u1_u1_7717_wire <= (zero_result_7654 or div_by_0_trap_7595);
    -- flow through binary operator OR_u1_u1_7736_inst
    OR_u1_u1_7736_wire <= (EQ_u33_u1_7730_wire or EQ_u33_u1_7735_wire);
    -- flow through binary operator OR_u64_u64_7697_inst
    OR_u64_u64_7697_wire <= (MUX_7690_wire or MUX_7696_wire);
    -- flow through binary operator OR_u64_u64_7702_inst
    no_trap_result_7703 <= (OR_u64_u64_7697_wire or MUX_7701_wire);
    -- flow through binary operator XOR_u1_u1_7708_inst
    XOR_u1_u1_7708_wire <= (sdividend_7600 xor sdivisor_7610);
    volatile_operator_twos_complement_64_6909: twos_complement_64_Volatile port map(A => dividend_64_7605, B => inverted_dividend_64_7613); 
    volatile_operator_twos_complement_32_6912: twos_complement_32_Volatile port map(A => divisor_buffer, B => inverted_divisor_7625); 
    volatile_operator_u_cmp_32_6917: u_cmp_32_Volatile port map(a => udividend_l_7641, b => udivisor_7633, l => l_7647, g => g_7647, e => e_7647); 
    -- shared call operator group (3) : call_stmt_7685_call 
    u64_true_divide_revised_call_group_3: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_7685_call_req_0;
      call_stmt_7685_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_7685_call_req_1;
      call_stmt_7685_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= run_true_divide_7680(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      u64_true_divide_revised_call_group_3_gI: SplitGuardInterface generic map(name => "u64_true_divide_revised_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= udividend_7622 & udivisor_7633;
      QUOTIENT_7685 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 96,
        owidth => 96,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => u64_true_divide_revised_call_reqs(0),
          ackR => u64_true_divide_revised_call_acks(0),
          dataR => u64_true_divide_revised_call_data(95 downto 0),
          tagR => u64_true_divide_revised_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => u64_true_divide_revised_return_acks(0), -- cross-over
          ackL => u64_true_divide_revised_return_reqs(0), -- cross-over
          dataL => u64_true_divide_revised_return_data(63 downto 0),
          tagL => u64_true_divide_revised_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    volatile_operator_twos_complement_64_6937: twos_complement_64_Volatile port map(A => no_trap_result_7703, B => inverted_no_trap_result_7713); 
    -- 
  end Block; -- data_path
  -- 
end i32_div_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity i32_mul_calculate_sign_correction_Volatile is -- 
  port ( -- 
    signed_mul : in  std_logic_vector(0 downto 0);
    A : in  std_logic_vector(31 downto 0);
    B : in  std_logic_vector(31 downto 0);
    sign_correction : out  std_logic_vector(31 downto 0)-- 
  );
  -- 
end entity i32_mul_calculate_sign_correction_Volatile;
architecture i32_mul_calculate_sign_correction_Volatile_arch of i32_mul_calculate_sign_correction_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(65-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal signed_mul_buffer :  std_logic_vector(0 downto 0);
  signal A_buffer :  std_logic_vector(31 downto 0);
  signal B_buffer :  std_logic_vector(31 downto 0);
  -- output port buffer signals
  signal sign_correction_buffer :  std_logic_vector(31 downto 0);
  -- volatile/operator module components. 
  component twos_complement_32_Volatile is -- 
    port ( -- 
      A : in  std_logic_vector(31 downto 0);
      B : out  std_logic_vector(31 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  signed_mul_buffer <= signed_mul;
  A_buffer <= A;
  B_buffer <= B;
  -- output handling  -------------------------------------------------------
  sign_correction <= sign_correction_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal MUX_7815_wire : std_logic_vector(31 downto 0);
    signal MUX_7819_wire : std_logic_vector(31 downto 0);
    signal OR_u1_u1_7828_wire : std_logic_vector(0 downto 0);
    signal X_7821 : std_logic_vector(31 downto 0);
    signal inverted_X_7824 : std_logic_vector(31 downto 0);
    signal konst_7803_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7808_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7814_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7818_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7830_wire_constant : std_logic_vector(31 downto 0);
    signal sA_7805 : std_logic_vector(0 downto 0);
    signal sB_7810 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_7803_wire_constant <= "00000000000000000000000000011111";
    konst_7808_wire_constant <= "00000000000000000000000000011111";
    konst_7814_wire_constant <= "00000000000000000000000000000000";
    konst_7818_wire_constant <= "00000000000000000000000000000000";
    konst_7830_wire_constant <= "00000000000000000000000000000000";
    -- flow-through select operator MUX_7815_inst
    MUX_7815_wire <= B_buffer when (sA_7805(0) /=  '0') else konst_7814_wire_constant;
    -- flow-through select operator MUX_7819_inst
    MUX_7819_wire <= A_buffer when (sB_7810(0) /=  '0') else konst_7818_wire_constant;
    -- flow-through select operator MUX_7831_inst
    sign_correction_buffer <= inverted_X_7824 when (OR_u1_u1_7828_wire(0) /=  '0') else konst_7830_wire_constant;
    -- flow through binary operator ADD_u32_u32_7820_inst
    X_7821 <= std_logic_vector(unsigned(MUX_7815_wire) + unsigned(MUX_7819_wire));
    -- flow through binary operator BITSEL_u32_u1_7804_inst
    process(A_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(A_buffer, konst_7803_wire_constant, tmp_var);
      sA_7805 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_7809_inst
    process(B_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(B_buffer, konst_7808_wire_constant, tmp_var);
      sB_7810 <= tmp_var; --
    end process;
    -- flow through binary operator OR_u1_u1_7828_inst
    OR_u1_u1_7828_wire <= (sA_7805 or sB_7810);
    volatile_operator_twos_complement_32_7035: twos_complement_32_Volatile port map(A => X_7821, B => inverted_X_7824); 
    -- 
  end Block; -- data_path
  -- 
end i32_mul_calculate_sign_correction_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity i32_mulscc_Volatile is -- 
  port ( -- 
    y_in : in  std_logic_vector(31 downto 0);
    A : in  std_logic_vector(31 downto 0);
    B : in  std_logic_vector(31 downto 0);
    Ni : in  std_logic_vector(0 downto 0);
    Zi : in  std_logic_vector(0 downto 0);
    Vi : in  std_logic_vector(0 downto 0);
    Ci : in  std_logic_vector(0 downto 0);
    y_out : out  std_logic_vector(31 downto 0);
    result : out  std_logic_vector(31 downto 0);
    No : out  std_logic_vector(0 downto 0);
    Zo : out  std_logic_vector(0 downto 0);
    Vo : out  std_logic_vector(0 downto 0);
    Co : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity i32_mulscc_Volatile;
architecture i32_mulscc_Volatile_arch of i32_mulscc_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(100-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal y_in_buffer :  std_logic_vector(31 downto 0);
  signal A_buffer :  std_logic_vector(31 downto 0);
  signal B_buffer :  std_logic_vector(31 downto 0);
  signal Ni_buffer :  std_logic_vector(0 downto 0);
  signal Zi_buffer :  std_logic_vector(0 downto 0);
  signal Vi_buffer :  std_logic_vector(0 downto 0);
  signal Ci_buffer :  std_logic_vector(0 downto 0);
  -- output port buffer signals
  signal y_out_buffer :  std_logic_vector(31 downto 0);
  signal result_buffer :  std_logic_vector(31 downto 0);
  signal No_buffer :  std_logic_vector(0 downto 0);
  signal Zo_buffer :  std_logic_vector(0 downto 0);
  signal Vo_buffer :  std_logic_vector(0 downto 0);
  signal Co_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  component i32_add_sub_Volatile is -- 
    port ( -- 
      subtract_flag : in  std_logic_vector(0 downto 0);
      with_carry : in  std_logic_vector(0 downto 0);
      set_cc : in  std_logic_vector(0 downto 0);
      tagged_op : in  std_logic_vector(0 downto 0);
      trap_on_ovflow : in  std_logic_vector(0 downto 0);
      Ni : in  std_logic_vector(0 downto 0);
      Zi : in  std_logic_vector(0 downto 0);
      Vi : in  std_logic_vector(0 downto 0);
      Ci : in  std_logic_vector(0 downto 0);
      x : in  std_logic_vector(31 downto 0);
      y : in  std_logic_vector(31 downto 0);
      result : out  std_logic_vector(31 downto 0);
      No : out  std_logic_vector(0 downto 0);
      Zo : out  std_logic_vector(0 downto 0);
      Vo : out  std_logic_vector(0 downto 0);
      Co : out  std_logic_vector(0 downto 0);
      overflow_trap : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  y_in_buffer <= y_in;
  A_buffer <= A;
  B_buffer <= B;
  Ni_buffer <= Ni;
  Zi_buffer <= Zi;
  Vi_buffer <= Vi;
  Ci_buffer <= Ci;
  -- output handling  -------------------------------------------------------
  y_out <= y_out_buffer;
  result <= result_buffer;
  No <= No_buffer;
  Zo <= Zo_buffer;
  Vo <= Vo_buffer;
  Co <= Co_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_7977_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7980_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7985_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7987_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7993_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7999_wire : std_logic_vector(0 downto 0);
    signal Ap_7919 : std_logic_vector(31 downto 0);
    signal BITSEL_u32_u1_7928_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_7959_wire : std_logic_vector(0 downto 0);
    signal Bp_7932 : std_logic_vector(31 downto 0);
    signal NOT_u1_u1_7979_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_7982_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_7984_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_7995_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_7998_wire : std_logic_vector(0 downto 0);
    signal R_ZERO_1_7939_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_7940_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_7941_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_7942_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_7943_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_7944_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_7945_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_7946_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_32_7930_wire_constant : std_logic_vector(31 downto 0);
    signal XOR_u1_u1_7915_wire : std_logic_vector(0 downto 0);
    signal ignC_7955 : std_logic_vector(0 downto 0);
    signal ignN_7955 : std_logic_vector(0 downto 0);
    signal ignTrp_7955 : std_logic_vector(0 downto 0);
    signal ignV_7955 : std_logic_vector(0 downto 0);
    signal ignZ_7955 : std_logic_vector(0 downto 0);
    signal konst_7922_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7927_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7935_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7938_wire_constant : std_logic_vector(0 downto 0);
    signal konst_7958_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7966_wire_constant : std_logic_vector(31 downto 0);
    signal konst_7971_wire_constant : std_logic_vector(31 downto 0);
    signal raw_result_7955 : std_logic_vector(31 downto 0);
    signal sA_7924 : std_logic_vector(0 downto 0);
    signal sB_7937 : std_logic_vector(0 downto 0);
    signal slice_7917_wire : std_logic_vector(30 downto 0);
    signal slice_7961_wire : std_logic_vector(30 downto 0);
    -- 
  begin -- 
    R_ZERO_1_7939_wire_constant <= "0";
    R_ZERO_1_7940_wire_constant <= "0";
    R_ZERO_1_7941_wire_constant <= "0";
    R_ZERO_1_7942_wire_constant <= "0";
    R_ZERO_1_7943_wire_constant <= "0";
    R_ZERO_1_7944_wire_constant <= "0";
    R_ZERO_1_7945_wire_constant <= "0";
    R_ZERO_1_7946_wire_constant <= "0";
    R_ZERO_32_7930_wire_constant <= "00000000000000000000000000000000";
    konst_7922_wire_constant <= "00000000000000000000000000011111";
    konst_7927_wire_constant <= "00000000000000000000000000000000";
    konst_7935_wire_constant <= "00000000000000000000000000011111";
    konst_7938_wire_constant <= "0";
    konst_7958_wire_constant <= "00000000000000000000000000000000";
    konst_7966_wire_constant <= "00000000000000000000000000011111";
    konst_7971_wire_constant <= "00000000000000000000000000000000";
    -- flow-through select operator MUX_7931_inst
    Bp_7932 <= B_buffer when (BITSEL_u32_u1_7928_wire(0) /=  '0') else R_ZERO_32_7930_wire_constant;
    -- flow-through slice operator slice_7917_inst
    slice_7917_wire <= A_buffer(31 downto 1);
    -- flow-through slice operator slice_7961_inst
    slice_7961_wire <= y_in_buffer(31 downto 1);
    -- interlock W_result_8002_inst
    process(raw_result_7955) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := raw_result_7955(31 downto 0);
      result_buffer <= tmp_var; -- 
    end process;
    -- flow through binary operator AND_u1_u1_7977_inst
    AND_u1_u1_7977_wire <= (sA_7924 and sB_7937);
    -- flow through binary operator AND_u1_u1_7980_inst
    AND_u1_u1_7980_wire <= (AND_u1_u1_7977_wire and NOT_u1_u1_7979_wire);
    -- flow through binary operator AND_u1_u1_7985_inst
    AND_u1_u1_7985_wire <= (NOT_u1_u1_7982_wire and NOT_u1_u1_7984_wire);
    -- flow through binary operator AND_u1_u1_7987_inst
    AND_u1_u1_7987_wire <= (AND_u1_u1_7985_wire and No_buffer);
    -- flow through binary operator AND_u1_u1_7993_inst
    AND_u1_u1_7993_wire <= (sA_7924 and sB_7937);
    -- flow through binary operator AND_u1_u1_7999_inst
    AND_u1_u1_7999_wire <= (NOT_u1_u1_7995_wire and OR_u1_u1_7998_wire);
    -- flow through binary operator BITSEL_u32_u1_7923_inst
    process(Ap_7919) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(Ap_7919, konst_7922_wire_constant, tmp_var);
      sA_7924 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_7928_inst
    process(y_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(y_in_buffer, konst_7927_wire_constant, tmp_var);
      BITSEL_u32_u1_7928_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_7936_inst
    process(Bp_7932) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(Bp_7932, konst_7935_wire_constant, tmp_var);
      sB_7937 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_7959_inst
    process(A_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(A_buffer, konst_7958_wire_constant, tmp_var);
      BITSEL_u32_u1_7959_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_7967_inst
    process(raw_result_7955) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(raw_result_7955, konst_7966_wire_constant, tmp_var);
      No_buffer <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u32_7918_inst
    process(XOR_u1_u1_7915_wire, slice_7917_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(XOR_u1_u1_7915_wire, slice_7917_wire, tmp_var);
      Ap_7919 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u32_7962_inst
    process(BITSEL_u32_u1_7959_wire, slice_7961_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(BITSEL_u32_u1_7959_wire, slice_7961_wire, tmp_var);
      y_out_buffer <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_7972_inst
    process(raw_result_7955) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(raw_result_7955, konst_7971_wire_constant, tmp_var);
      Zo_buffer <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_7979_inst
    process(No_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", No_buffer, tmp_var);
      NOT_u1_u1_7979_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_7982_inst
    process(sA_7924) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", sA_7924, tmp_var);
      NOT_u1_u1_7982_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_7984_inst
    process(sB_7937) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", sB_7937, tmp_var);
      NOT_u1_u1_7984_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_7995_inst
    process(No_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", No_buffer, tmp_var);
      NOT_u1_u1_7995_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_7988_inst
    Vo_buffer <= (AND_u1_u1_7980_wire or AND_u1_u1_7987_wire);
    -- flow through binary operator OR_u1_u1_7998_inst
    OR_u1_u1_7998_wire <= (sA_7924 or sB_7937);
    -- flow through binary operator OR_u1_u1_8000_inst
    Co_buffer <= (AND_u1_u1_7993_wire or AND_u1_u1_7999_wire);
    -- flow through binary operator XOR_u1_u1_7915_inst
    XOR_u1_u1_7915_wire <= (Ni_buffer xor Vi_buffer);
    volatile_operator_i32_add_sub_7281: i32_add_sub_Volatile port map(subtract_flag => konst_7938_wire_constant, with_carry => R_ZERO_1_7939_wire_constant, set_cc => R_ZERO_1_7940_wire_constant, tagged_op => R_ZERO_1_7941_wire_constant, trap_on_ovflow => R_ZERO_1_7942_wire_constant, Ni => R_ZERO_1_7943_wire_constant, Zi => R_ZERO_1_7944_wire_constant, Vi => R_ZERO_1_7945_wire_constant, Ci => R_ZERO_1_7946_wire_constant, x => Ap_7919, y => Bp_7932, result => raw_result_7955, No => ignN_7955, Zo => ignZ_7955, Vo => ignV_7955, Co => ignC_7955, overflow_trap => ignTrp_7955); 
    -- 
  end Block; -- data_path
  -- 
end i32_mulscc_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity i32_shift_Volatile is -- 
  port ( -- 
    is_sll : in  std_logic_vector(0 downto 0);
    is_srl : in  std_logic_vector(0 downto 0);
    is_sra : in  std_logic_vector(0 downto 0);
    x : in  std_logic_vector(31 downto 0);
    shift_amount : in  std_logic_vector(31 downto 0);
    result : out  std_logic_vector(31 downto 0)-- 
  );
  -- 
end entity i32_shift_Volatile;
architecture i32_shift_Volatile_arch of i32_shift_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(67-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal is_sll_buffer :  std_logic_vector(0 downto 0);
  signal is_srl_buffer :  std_logic_vector(0 downto 0);
  signal is_sra_buffer :  std_logic_vector(0 downto 0);
  signal x_buffer :  std_logic_vector(31 downto 0);
  signal shift_amount_buffer :  std_logic_vector(31 downto 0);
  -- output port buffer signals
  signal result_buffer :  std_logic_vector(31 downto 0);
  -- volatile/operator module components. 
  component i32_sll_Volatile is -- 
    port ( -- 
      X : in  std_logic_vector(31 downto 0);
      S : in  std_logic_vector(4 downto 0);
      Y : out  std_logic_vector(31 downto 0)-- 
    );
    -- 
  end component; 
  component i32_srl_Volatile is -- 
    port ( -- 
      X : in  std_logic_vector(31 downto 0);
      S : in  std_logic_vector(4 downto 0);
      Y : out  std_logic_vector(31 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  is_sll_buffer <= is_sll;
  is_srl_buffer <= is_srl;
  is_sra_buffer <= is_sra;
  x_buffer <= x;
  shift_amount_buffer <= shift_amount;
  -- output handling  -------------------------------------------------------
  result <= result_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_8213_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_8209_wire : std_logic_vector(0 downto 0);
    signal MUX_8237_wire : std_logic_vector(31 downto 0);
    signal MUX_8241_wire : std_logic_vector(31 downto 0);
    signal MUX_8246_wire : std_logic_vector(31 downto 0);
    signal NEQ_u5_u1_8212_wire : std_logic_vector(0 downto 0);
    signal NOT_u32_u32_8186_wire_constant : std_logic_vector(31 downto 0);
    signal OR_u32_u32_8242_wire : std_logic_vector(31 downto 0);
    signal R_ZERO_32_8215_wire_constant : std_logic_vector(31 downto 0);
    signal S6_8177 : std_logic_vector(5 downto 0);
    signal SUB_u6_u6_8194_wire : std_logic_vector(5 downto 0);
    signal S_8181 : std_logic_vector(4 downto 0);
    signal konst_8192_wire_constant : std_logic_vector(5 downto 0);
    signal konst_8208_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8211_wire_constant : std_logic_vector(4 downto 0);
    signal konst_8236_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8240_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8245_wire_constant : std_logic_vector(31 downto 0);
    signal result_sll_8201 : std_logic_vector(31 downto 0);
    signal result_sra_8222 : std_logic_vector(31 downto 0);
    signal result_srl_8205 : std_logic_vector(31 downto 0);
    signal slice_8195_wire : std_logic_vector(4 downto 0);
    signal sll_S_8197 : std_logic_vector(4 downto 0);
    signal sll_X_8188 : std_logic_vector(31 downto 0);
    signal sra_mask_8217 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    NOT_u32_u32_8186_wire_constant <= "11111111111111111111111111111111";
    R_ZERO_32_8215_wire_constant <= "00000000000000000000000000000000";
    konst_8192_wire_constant <= "100000";
    konst_8208_wire_constant <= "00000000000000000000000000011111";
    konst_8211_wire_constant <= "00000";
    konst_8236_wire_constant <= "00000000000000000000000000000000";
    konst_8240_wire_constant <= "00000000000000000000000000000000";
    konst_8245_wire_constant <= "00000000000000000000000000000000";
    -- flow-through select operator MUX_8187_inst
    sll_X_8188 <= x_buffer when (is_sll_buffer(0) /=  '0') else NOT_u32_u32_8186_wire_constant;
    -- flow-through select operator MUX_8196_inst
    sll_S_8197 <= S_8181 when (is_sll_buffer(0) /=  '0') else slice_8195_wire;
    -- flow-through select operator MUX_8216_inst
    sra_mask_8217 <= result_sll_8201 when (AND_u1_u1_8213_wire(0) /=  '0') else R_ZERO_32_8215_wire_constant;
    -- flow-through select operator MUX_8237_inst
    MUX_8237_wire <= result_sll_8201 when (is_sll_buffer(0) /=  '0') else konst_8236_wire_constant;
    -- flow-through select operator MUX_8241_inst
    MUX_8241_wire <= result_srl_8205 when (is_srl_buffer(0) /=  '0') else konst_8240_wire_constant;
    -- flow-through select operator MUX_8246_inst
    MUX_8246_wire <= result_sra_8222 when (is_sra_buffer(0) /=  '0') else konst_8245_wire_constant;
    -- flow-through slice operator slice_8176_inst
    S6_8177 <= shift_amount_buffer(5 downto 0);
    -- flow-through slice operator slice_8180_inst
    S_8181 <= shift_amount_buffer(4 downto 0);
    -- flow-through slice operator slice_8195_inst
    slice_8195_wire <= SUB_u6_u6_8194_wire(4 downto 0);
    -- flow through binary operator AND_u1_u1_8213_inst
    AND_u1_u1_8213_wire <= (BITSEL_u32_u1_8209_wire and NEQ_u5_u1_8212_wire);
    -- flow through binary operator BITSEL_u32_u1_8209_inst
    process(x_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(x_buffer, konst_8208_wire_constant, tmp_var);
      BITSEL_u32_u1_8209_wire <= tmp_var; --
    end process;
    -- flow through binary operator NEQ_u5_u1_8212_inst
    process(S_8181) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(S_8181, konst_8211_wire_constant, tmp_var);
      NEQ_u5_u1_8212_wire <= tmp_var; --
    end process;
    -- flow through binary operator OR_u32_u32_8221_inst
    result_sra_8222 <= (result_srl_8205 or sra_mask_8217);
    -- flow through binary operator OR_u32_u32_8242_inst
    OR_u32_u32_8242_wire <= (MUX_8237_wire or MUX_8241_wire);
    -- flow through binary operator OR_u32_u32_8247_inst
    result_buffer <= (OR_u32_u32_8242_wire or MUX_8246_wire);
    -- flow through binary operator SUB_u6_u6_8194_inst
    SUB_u6_u6_8194_wire <= std_logic_vector(unsigned(konst_8192_wire_constant) - unsigned(S6_8177));
    volatile_operator_i32_sll_7543: i32_sll_Volatile port map(X => sll_X_8188, S => sll_S_8197, Y => result_sll_8201); 
    volatile_operator_i32_srl_7544: i32_srl_Volatile port map(X => x_buffer, S => S_8181, Y => result_srl_8205); 
    -- 
  end Block; -- data_path
  -- 
end i32_shift_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity i32_sll_Volatile is -- 
  port ( -- 
    X : in  std_logic_vector(31 downto 0);
    S : in  std_logic_vector(4 downto 0);
    Y : out  std_logic_vector(31 downto 0)-- 
  );
  -- 
end entity i32_sll_Volatile;
architecture i32_sll_Volatile_arch of i32_sll_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(37-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal X_buffer :  std_logic_vector(31 downto 0);
  signal S_buffer :  std_logic_vector(4 downto 0);
  -- output port buffer signals
  signal Y_buffer :  std_logic_vector(31 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  X_buffer <= X;
  S_buffer <= S;
  -- output handling  -------------------------------------------------------
  Y <= Y_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u5_u1_8054_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u5_u1_8065_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u5_u1_8076_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u5_u1_8087_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u5_u1_8098_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u16_u32_8102_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u24_u32_8091_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u28_u32_8080_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u30_u32_8069_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u31_u32_8058_wire : std_logic_vector(31 downto 0);
    signal R_ZERO_16_8101_wire_constant : std_logic_vector(15 downto 0);
    signal R_ZERO_1_8057_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_2_8068_wire_constant : std_logic_vector(1 downto 0);
    signal R_ZERO_4_8079_wire_constant : std_logic_vector(3 downto 0);
    signal R_ZERO_8_8090_wire_constant : std_logic_vector(7 downto 0);
    signal X0_8061 : std_logic_vector(31 downto 0);
    signal X1_8072 : std_logic_vector(31 downto 0);
    signal X2_8083 : std_logic_vector(31 downto 0);
    signal X3_8094 : std_logic_vector(31 downto 0);
    signal konst_8053_wire_constant : std_logic_vector(4 downto 0);
    signal konst_8064_wire_constant : std_logic_vector(4 downto 0);
    signal konst_8075_wire_constant : std_logic_vector(4 downto 0);
    signal konst_8086_wire_constant : std_logic_vector(4 downto 0);
    signal konst_8097_wire_constant : std_logic_vector(4 downto 0);
    signal slice_8056_wire : std_logic_vector(30 downto 0);
    signal slice_8067_wire : std_logic_vector(29 downto 0);
    signal slice_8078_wire : std_logic_vector(27 downto 0);
    signal slice_8089_wire : std_logic_vector(23 downto 0);
    signal slice_8100_wire : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ZERO_16_8101_wire_constant <= "0000000000000000";
    R_ZERO_1_8057_wire_constant <= "0";
    R_ZERO_2_8068_wire_constant <= "00";
    R_ZERO_4_8079_wire_constant <= "0000";
    R_ZERO_8_8090_wire_constant <= "00000000";
    konst_8053_wire_constant <= "00000";
    konst_8064_wire_constant <= "00001";
    konst_8075_wire_constant <= "00010";
    konst_8086_wire_constant <= "00011";
    konst_8097_wire_constant <= "00100";
    -- flow-through select operator MUX_8060_inst
    X0_8061 <= CONCAT_u31_u32_8058_wire when (BITSEL_u5_u1_8054_wire(0) /=  '0') else X_buffer;
    -- flow-through select operator MUX_8071_inst
    X1_8072 <= CONCAT_u30_u32_8069_wire when (BITSEL_u5_u1_8065_wire(0) /=  '0') else X0_8061;
    -- flow-through select operator MUX_8082_inst
    X2_8083 <= CONCAT_u28_u32_8080_wire when (BITSEL_u5_u1_8076_wire(0) /=  '0') else X1_8072;
    -- flow-through select operator MUX_8093_inst
    X3_8094 <= CONCAT_u24_u32_8091_wire when (BITSEL_u5_u1_8087_wire(0) /=  '0') else X2_8083;
    -- flow-through select operator MUX_8104_inst
    Y_buffer <= CONCAT_u16_u32_8102_wire when (BITSEL_u5_u1_8098_wire(0) /=  '0') else X3_8094;
    -- flow-through slice operator slice_8056_inst
    slice_8056_wire <= X_buffer(30 downto 0);
    -- flow-through slice operator slice_8067_inst
    slice_8067_wire <= X0_8061(29 downto 0);
    -- flow-through slice operator slice_8078_inst
    slice_8078_wire <= X1_8072(27 downto 0);
    -- flow-through slice operator slice_8089_inst
    slice_8089_wire <= X2_8083(23 downto 0);
    -- flow-through slice operator slice_8100_inst
    slice_8100_wire <= X3_8094(15 downto 0);
    -- flow through binary operator BITSEL_u5_u1_8054_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_8053_wire_constant, tmp_var);
      BITSEL_u5_u1_8054_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u5_u1_8065_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_8064_wire_constant, tmp_var);
      BITSEL_u5_u1_8065_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u5_u1_8076_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_8075_wire_constant, tmp_var);
      BITSEL_u5_u1_8076_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u5_u1_8087_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_8086_wire_constant, tmp_var);
      BITSEL_u5_u1_8087_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u5_u1_8098_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_8097_wire_constant, tmp_var);
      BITSEL_u5_u1_8098_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u16_u32_8102_inst
    process(slice_8100_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_8100_wire, R_ZERO_16_8101_wire_constant, tmp_var);
      CONCAT_u16_u32_8102_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u24_u32_8091_inst
    process(slice_8089_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_8089_wire, R_ZERO_8_8090_wire_constant, tmp_var);
      CONCAT_u24_u32_8091_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u28_u32_8080_inst
    process(slice_8078_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_8078_wire, R_ZERO_4_8079_wire_constant, tmp_var);
      CONCAT_u28_u32_8080_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u30_u32_8069_inst
    process(slice_8067_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_8067_wire, R_ZERO_2_8068_wire_constant, tmp_var);
      CONCAT_u30_u32_8069_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u31_u32_8058_inst
    process(slice_8056_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_8056_wire, R_ZERO_1_8057_wire_constant, tmp_var);
      CONCAT_u31_u32_8058_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end i32_sll_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity i32_srl_Volatile is -- 
  port ( -- 
    X : in  std_logic_vector(31 downto 0);
    S : in  std_logic_vector(4 downto 0);
    Y : out  std_logic_vector(31 downto 0)-- 
  );
  -- 
end entity i32_srl_Volatile;
architecture i32_srl_Volatile_arch of i32_srl_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(37-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal X_buffer :  std_logic_vector(31 downto 0);
  signal S_buffer :  std_logic_vector(4 downto 0);
  -- output port buffer signals
  signal Y_buffer :  std_logic_vector(31 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  X_buffer <= X;
  S_buffer <= S;
  -- output handling  -------------------------------------------------------
  Y <= Y_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u5_u1_8114_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u5_u1_8125_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u5_u1_8136_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u5_u1_8147_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u5_u1_8158_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u16_u32_8162_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u1_u32_8118_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u2_u32_8129_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u4_u32_8140_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u8_u32_8151_wire : std_logic_vector(31 downto 0);
    signal R_ZERO_16_8159_wire_constant : std_logic_vector(15 downto 0);
    signal R_ZERO_1_8115_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_2_8126_wire_constant : std_logic_vector(1 downto 0);
    signal R_ZERO_4_8137_wire_constant : std_logic_vector(3 downto 0);
    signal R_ZERO_8_8148_wire_constant : std_logic_vector(7 downto 0);
    signal X0_8121 : std_logic_vector(31 downto 0);
    signal X1_8132 : std_logic_vector(31 downto 0);
    signal X2_8143 : std_logic_vector(31 downto 0);
    signal X3_8154 : std_logic_vector(31 downto 0);
    signal konst_8113_wire_constant : std_logic_vector(4 downto 0);
    signal konst_8124_wire_constant : std_logic_vector(4 downto 0);
    signal konst_8135_wire_constant : std_logic_vector(4 downto 0);
    signal konst_8146_wire_constant : std_logic_vector(4 downto 0);
    signal konst_8157_wire_constant : std_logic_vector(4 downto 0);
    signal slice_8117_wire : std_logic_vector(30 downto 0);
    signal slice_8128_wire : std_logic_vector(29 downto 0);
    signal slice_8139_wire : std_logic_vector(27 downto 0);
    signal slice_8150_wire : std_logic_vector(23 downto 0);
    signal slice_8161_wire : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ZERO_16_8159_wire_constant <= "0000000000000000";
    R_ZERO_1_8115_wire_constant <= "0";
    R_ZERO_2_8126_wire_constant <= "00";
    R_ZERO_4_8137_wire_constant <= "0000";
    R_ZERO_8_8148_wire_constant <= "00000000";
    konst_8113_wire_constant <= "00000";
    konst_8124_wire_constant <= "00001";
    konst_8135_wire_constant <= "00010";
    konst_8146_wire_constant <= "00011";
    konst_8157_wire_constant <= "00100";
    -- flow-through select operator MUX_8120_inst
    X0_8121 <= CONCAT_u1_u32_8118_wire when (BITSEL_u5_u1_8114_wire(0) /=  '0') else X_buffer;
    -- flow-through select operator MUX_8131_inst
    X1_8132 <= CONCAT_u2_u32_8129_wire when (BITSEL_u5_u1_8125_wire(0) /=  '0') else X0_8121;
    -- flow-through select operator MUX_8142_inst
    X2_8143 <= CONCAT_u4_u32_8140_wire when (BITSEL_u5_u1_8136_wire(0) /=  '0') else X1_8132;
    -- flow-through select operator MUX_8153_inst
    X3_8154 <= CONCAT_u8_u32_8151_wire when (BITSEL_u5_u1_8147_wire(0) /=  '0') else X2_8143;
    -- flow-through select operator MUX_8164_inst
    Y_buffer <= CONCAT_u16_u32_8162_wire when (BITSEL_u5_u1_8158_wire(0) /=  '0') else X3_8154;
    -- flow-through slice operator slice_8117_inst
    slice_8117_wire <= X_buffer(31 downto 1);
    -- flow-through slice operator slice_8128_inst
    slice_8128_wire <= X0_8121(31 downto 2);
    -- flow-through slice operator slice_8139_inst
    slice_8139_wire <= X1_8132(31 downto 4);
    -- flow-through slice operator slice_8150_inst
    slice_8150_wire <= X2_8143(31 downto 8);
    -- flow-through slice operator slice_8161_inst
    slice_8161_wire <= X3_8154(31 downto 16);
    -- flow through binary operator BITSEL_u5_u1_8114_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_8113_wire_constant, tmp_var);
      BITSEL_u5_u1_8114_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u5_u1_8125_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_8124_wire_constant, tmp_var);
      BITSEL_u5_u1_8125_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u5_u1_8136_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_8135_wire_constant, tmp_var);
      BITSEL_u5_u1_8136_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u5_u1_8147_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_8146_wire_constant, tmp_var);
      BITSEL_u5_u1_8147_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u5_u1_8158_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_8157_wire_constant, tmp_var);
      BITSEL_u5_u1_8158_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u16_u32_8162_inst
    process(R_ZERO_16_8159_wire_constant, slice_8161_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_16_8159_wire_constant, slice_8161_wire, tmp_var);
      CONCAT_u16_u32_8162_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u32_8118_inst
    process(R_ZERO_1_8115_wire_constant, slice_8117_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_1_8115_wire_constant, slice_8117_wire, tmp_var);
      CONCAT_u1_u32_8118_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u32_8129_inst
    process(R_ZERO_2_8126_wire_constant, slice_8128_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_2_8126_wire_constant, slice_8128_wire, tmp_var);
      CONCAT_u2_u32_8129_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u4_u32_8140_inst
    process(R_ZERO_4_8137_wire_constant, slice_8139_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_4_8137_wire_constant, slice_8139_wire, tmp_var);
      CONCAT_u4_u32_8140_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u8_u32_8151_inst
    process(R_ZERO_8_8148_wire_constant, slice_8150_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_8_8148_wire_constant, slice_8150_wire, tmp_var);
      CONCAT_u8_u32_8151_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end i32_srl_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity increment_16_Volatile is -- 
  port ( -- 
    A : in  std_logic_vector(15 downto 0);
    B : out  std_logic_vector(15 downto 0)-- 
  );
  -- 
end entity increment_16_Volatile;
architecture increment_16_Volatile_arch of increment_16_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(16-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal A_buffer :  std_logic_vector(15 downto 0);
  -- output port buffer signals
  signal B_buffer :  std_logic_vector(15 downto 0);
  -- volatile/operator module components. 
  component increment_8_Volatile is -- 
    port ( -- 
      cA : in  std_logic_vector(7 downto 0);
      B : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  A_buffer <= A;
  -- output handling  -------------------------------------------------------
  B <= B_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AH_7194 : std_logic_vector(7 downto 0);
    signal AL_7198 : std_logic_vector(7 downto 0);
    signal BL_7201 : std_logic_vector(7 downto 0);
    signal EQ_u8_u1_7209_wire : std_logic_vector(0 downto 0);
    signal MUX_7212_wire : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_7207_wire : std_logic_vector(7 downto 0);
    signal konst_7208_wire_constant : std_logic_vector(7 downto 0);
    signal tBH_7204 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_7208_wire_constant <= "00000000";
    -- flow-through select operator MUX_7212_inst
    MUX_7212_wire <= tBH_7204 when (EQ_u8_u1_7209_wire(0) /=  '0') else AH_7194;
    -- flow-through slice operator slice_7193_inst
    AH_7194 <= A_buffer(15 downto 8);
    -- flow-through slice operator slice_7197_inst
    AL_7198 <= A_buffer(7 downto 0);
    -- flow through binary operator CONCAT_u8_u16_7214_inst
    process(MUX_7212_wire, BL_7201) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_7212_wire, BL_7201, tmp_var);
      B_buffer <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u8_u1_7209_inst
    process(NOT_u8_u8_7207_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(NOT_u8_u8_7207_wire, konst_7208_wire_constant, tmp_var);
      EQ_u8_u1_7209_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u8_u8_7207_inst
    process(AL_7198) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", AL_7198, tmp_var);
      NOT_u8_u8_7207_wire <= tmp_var; -- 
    end process;
    volatile_operator_increment_8_6031: increment_8_Volatile port map(cA => AL_7198, B => BL_7201); 
    volatile_operator_increment_8_6032: increment_8_Volatile port map(cA => AH_7194, B => tBH_7204); 
    -- 
  end Block; -- data_path
  -- 
end increment_16_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity increment_32_Volatile is -- 
  port ( -- 
    A : in  std_logic_vector(31 downto 0);
    B : out  std_logic_vector(31 downto 0)-- 
  );
  -- 
end entity increment_32_Volatile;
architecture increment_32_Volatile_arch of increment_32_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(32-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal A_buffer :  std_logic_vector(31 downto 0);
  -- output port buffer signals
  signal B_buffer :  std_logic_vector(31 downto 0);
  -- volatile/operator module components. 
  component increment_16_Volatile is -- 
    port ( -- 
      A : in  std_logic_vector(15 downto 0);
      B : out  std_logic_vector(15 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  A_buffer <= A;
  -- output handling  -------------------------------------------------------
  B <= B_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AH_7223 : std_logic_vector(15 downto 0);
    signal AL_7227 : std_logic_vector(15 downto 0);
    signal BL_7230 : std_logic_vector(15 downto 0);
    signal EQ_u16_u1_7238_wire : std_logic_vector(0 downto 0);
    signal MUX_7241_wire : std_logic_vector(15 downto 0);
    signal NOT_u16_u16_7236_wire : std_logic_vector(15 downto 0);
    signal konst_7237_wire_constant : std_logic_vector(15 downto 0);
    signal tBH_7233 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    konst_7237_wire_constant <= "0000000000000000";
    -- flow-through select operator MUX_7241_inst
    MUX_7241_wire <= tBH_7233 when (EQ_u16_u1_7238_wire(0) /=  '0') else AH_7223;
    -- flow-through slice operator slice_7222_inst
    AH_7223 <= A_buffer(31 downto 16);
    -- flow-through slice operator slice_7226_inst
    AL_7227 <= A_buffer(15 downto 0);
    -- flow through binary operator CONCAT_u16_u32_7243_inst
    process(MUX_7241_wire, BL_7230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_7241_wire, BL_7230, tmp_var);
      B_buffer <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u16_u1_7238_inst
    process(NOT_u16_u16_7236_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(NOT_u16_u16_7236_wire, konst_7237_wire_constant, tmp_var);
      EQ_u16_u1_7238_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u16_u16_7236_inst
    process(AL_7227) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", AL_7227, tmp_var);
      NOT_u16_u16_7236_wire <= tmp_var; -- 
    end process;
    volatile_operator_increment_16_6055: increment_16_Volatile port map(A => AL_7227, B => BL_7230); 
    volatile_operator_increment_16_6056: increment_16_Volatile port map(A => AH_7223, B => tBH_7233); 
    -- 
  end Block; -- data_path
  -- 
end increment_32_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity increment_64_Volatile is -- 
  port ( -- 
    A : in  std_logic_vector(63 downto 0);
    B : out  std_logic_vector(63 downto 0)-- 
  );
  -- 
end entity increment_64_Volatile;
architecture increment_64_Volatile_arch of increment_64_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(64-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal A_buffer :  std_logic_vector(63 downto 0);
  -- output port buffer signals
  signal B_buffer :  std_logic_vector(63 downto 0);
  -- volatile/operator module components. 
  component increment_32_Volatile is -- 
    port ( -- 
      A : in  std_logic_vector(31 downto 0);
      B : out  std_logic_vector(31 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  A_buffer <= A;
  -- output handling  -------------------------------------------------------
  B <= B_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AH_7252 : std_logic_vector(31 downto 0);
    signal AL_7256 : std_logic_vector(31 downto 0);
    signal BL_7259 : std_logic_vector(31 downto 0);
    signal EQ_u32_u1_7267_wire : std_logic_vector(0 downto 0);
    signal MUX_7270_wire : std_logic_vector(31 downto 0);
    signal NOT_u32_u32_7265_wire : std_logic_vector(31 downto 0);
    signal konst_7266_wire_constant : std_logic_vector(31 downto 0);
    signal tBH_7262 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_7266_wire_constant <= "00000000000000000000000000000000";
    -- flow-through select operator MUX_7270_inst
    MUX_7270_wire <= tBH_7262 when (EQ_u32_u1_7267_wire(0) /=  '0') else AH_7252;
    -- flow-through slice operator slice_7251_inst
    AH_7252 <= A_buffer(63 downto 32);
    -- flow-through slice operator slice_7255_inst
    AL_7256 <= A_buffer(31 downto 0);
    -- flow through binary operator CONCAT_u32_u64_7272_inst
    process(MUX_7270_wire, BL_7259) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_7270_wire, BL_7259, tmp_var);
      B_buffer <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_7267_inst
    process(NOT_u32_u32_7265_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(NOT_u32_u32_7265_wire, konst_7266_wire_constant, tmp_var);
      EQ_u32_u1_7267_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u32_u32_7265_inst
    process(AL_7256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", AL_7256, tmp_var);
      NOT_u32_u32_7265_wire <= tmp_var; -- 
    end process;
    volatile_operator_increment_32_6079: increment_32_Volatile port map(A => AL_7256, B => BL_7259); 
    volatile_operator_increment_32_6080: increment_32_Volatile port map(A => AH_7252, B => tBH_7262); 
    -- 
  end Block; -- data_path
  -- 
end increment_64_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity increment_8_Volatile is -- 
  port ( -- 
    cA : in  std_logic_vector(7 downto 0);
    B : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity increment_8_Volatile;
architecture increment_8_Volatile_arch of increment_8_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal cA_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal B_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  cA_buffer <= cA;
  -- output handling  -------------------------------------------------------
  B <= B_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_7113_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7120_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7123_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7129_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7131_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7134_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7140_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7142_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7145_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7147_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7153_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7156_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7157_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7160_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7162_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u1_u2_7168_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_7171_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_7175_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_7178_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u4_7172_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_7179_wire : std_logic_vector(3 downto 0);
    signal b0_7098 : std_logic_vector(0 downto 0);
    signal b1_7094 : std_logic_vector(0 downto 0);
    signal b2_7090 : std_logic_vector(0 downto 0);
    signal b3_7086 : std_logic_vector(0 downto 0);
    signal b4_7082 : std_logic_vector(0 downto 0);
    signal b5_7078 : std_logic_vector(0 downto 0);
    signal b6_7074 : std_logic_vector(0 downto 0);
    signal c0_7101 : std_logic_vector(0 downto 0);
    signal c1_7104 : std_logic_vector(0 downto 0);
    signal c2_7109 : std_logic_vector(0 downto 0);
    signal c3_7116 : std_logic_vector(0 downto 0);
    signal c4_7125 : std_logic_vector(0 downto 0);
    signal c5_7136 : std_logic_vector(0 downto 0);
    signal c6_7149 : std_logic_vector(0 downto 0);
    signal c7_7164 : std_logic_vector(0 downto 0);
    signal c_7181 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    c0_7101 <= "1";
    -- flow-through slice operator slice_7073_inst
    b6_7074 <= cA_buffer(6 downto 6);
    -- flow-through slice operator slice_7077_inst
    b5_7078 <= cA_buffer(5 downto 5);
    -- flow-through slice operator slice_7081_inst
    b4_7082 <= cA_buffer(4 downto 4);
    -- flow-through slice operator slice_7085_inst
    b3_7086 <= cA_buffer(3 downto 3);
    -- flow-through slice operator slice_7089_inst
    b2_7090 <= cA_buffer(2 downto 2);
    -- flow-through slice operator slice_7093_inst
    b1_7094 <= cA_buffer(1 downto 1);
    -- flow-through slice operator slice_7097_inst
    b0_7098 <= cA_buffer(0 downto 0);
    -- interlock W_c1_7102_inst
    process(b0_7098) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := b0_7098(0 downto 0);
      c1_7104 <= tmp_var; -- 
    end process;
    -- flow through binary operator AND_u1_u1_7108_inst
    c2_7109 <= (b1_7094 and b0_7098);
    -- flow through binary operator AND_u1_u1_7113_inst
    AND_u1_u1_7113_wire <= (b2_7090 and b1_7094);
    -- flow through binary operator AND_u1_u1_7115_inst
    c3_7116 <= (AND_u1_u1_7113_wire and b0_7098);
    -- flow through binary operator AND_u1_u1_7120_inst
    AND_u1_u1_7120_wire <= (b3_7086 and b2_7090);
    -- flow through binary operator AND_u1_u1_7123_inst
    AND_u1_u1_7123_wire <= (b1_7094 and b0_7098);
    -- flow through binary operator AND_u1_u1_7124_inst
    c4_7125 <= (AND_u1_u1_7120_wire and AND_u1_u1_7123_wire);
    -- flow through binary operator AND_u1_u1_7129_inst
    AND_u1_u1_7129_wire <= (b4_7082 and b3_7086);
    -- flow through binary operator AND_u1_u1_7131_inst
    AND_u1_u1_7131_wire <= (AND_u1_u1_7129_wire and b2_7090);
    -- flow through binary operator AND_u1_u1_7134_inst
    AND_u1_u1_7134_wire <= (b1_7094 and b0_7098);
    -- flow through binary operator AND_u1_u1_7135_inst
    c5_7136 <= (AND_u1_u1_7131_wire and AND_u1_u1_7134_wire);
    -- flow through binary operator AND_u1_u1_7140_inst
    AND_u1_u1_7140_wire <= (b5_7078 and b4_7082);
    -- flow through binary operator AND_u1_u1_7142_inst
    AND_u1_u1_7142_wire <= (AND_u1_u1_7140_wire and b3_7086);
    -- flow through binary operator AND_u1_u1_7145_inst
    AND_u1_u1_7145_wire <= (b2_7090 and b1_7094);
    -- flow through binary operator AND_u1_u1_7147_inst
    AND_u1_u1_7147_wire <= (AND_u1_u1_7145_wire and b0_7098);
    -- flow through binary operator AND_u1_u1_7148_inst
    c6_7149 <= (AND_u1_u1_7142_wire and AND_u1_u1_7147_wire);
    -- flow through binary operator AND_u1_u1_7153_inst
    AND_u1_u1_7153_wire <= (b6_7074 and b5_7078);
    -- flow through binary operator AND_u1_u1_7156_inst
    AND_u1_u1_7156_wire <= (b4_7082 and b3_7086);
    -- flow through binary operator AND_u1_u1_7157_inst
    AND_u1_u1_7157_wire <= (AND_u1_u1_7153_wire and AND_u1_u1_7156_wire);
    -- flow through binary operator AND_u1_u1_7160_inst
    AND_u1_u1_7160_wire <= (b2_7090 and b1_7094);
    -- flow through binary operator AND_u1_u1_7162_inst
    AND_u1_u1_7162_wire <= (AND_u1_u1_7160_wire and b0_7098);
    -- flow through binary operator AND_u1_u1_7163_inst
    c7_7164 <= (AND_u1_u1_7157_wire and AND_u1_u1_7162_wire);
    -- flow through binary operator CONCAT_u1_u2_7168_inst
    process(c7_7164, c6_7149) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(c7_7164, c6_7149, tmp_var);
      CONCAT_u1_u2_7168_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_7171_inst
    process(c5_7136, c4_7125) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(c5_7136, c4_7125, tmp_var);
      CONCAT_u1_u2_7171_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_7175_inst
    process(c3_7116, c2_7109) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(c3_7116, c2_7109, tmp_var);
      CONCAT_u1_u2_7175_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_7178_inst
    process(c1_7104) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(c1_7104, c0_7101, tmp_var);
      CONCAT_u1_u2_7178_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u4_7172_inst
    process(CONCAT_u1_u2_7168_wire, CONCAT_u1_u2_7171_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_7168_wire, CONCAT_u1_u2_7171_wire, tmp_var);
      CONCAT_u2_u4_7172_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u4_7179_inst
    process(CONCAT_u1_u2_7175_wire, CONCAT_u1_u2_7178_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_7175_wire, CONCAT_u1_u2_7178_wire, tmp_var);
      CONCAT_u2_u4_7179_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u4_u8_7180_inst
    process(CONCAT_u2_u4_7172_wire, CONCAT_u2_u4_7179_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u4_7172_wire, CONCAT_u2_u4_7179_wire, tmp_var);
      c_7181 <= tmp_var; --
    end process;
    -- flow through binary operator XOR_u8_u8_7185_inst
    B_buffer <= (cA_buffer xor c_7181);
    -- 
  end Block; -- data_path
  -- 
end increment_8_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity iu_exec_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    iunit_register_file_read_access_response_pipe_read_req : out  std_logic_vector(0 downto 0);
    iunit_register_file_read_access_response_pipe_read_ack : in   std_logic_vector(0 downto 0);
    iunit_register_file_read_access_response_pipe_read_data : in   std_logic_vector(141 downto 0);
    teu_idispatch_to_iunit_exec_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_idispatch_to_iunit_exec_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_idispatch_to_iunit_exec_pipe_read_data : in   std_logic_vector(149 downto 0);
    noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_data : out  std_logic_vector(16 downto 0);
    noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_data : out  std_logic_vector(82 downto 0);
    noblock_iunit_exec_to_regfile_credit_return_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_iunit_exec_to_regfile_credit_return_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_iunit_exec_to_regfile_credit_return_pipe_write_data : out  std_logic_vector(0 downto 0);
    iunit_exec_fast_alu_result_to_writeback_pipe_write_req : out  std_logic_vector(0 downto 0);
    iunit_exec_fast_alu_result_to_writeback_pipe_write_ack : in   std_logic_vector(0 downto 0);
    iunit_exec_fast_alu_result_to_writeback_pipe_write_data : out  std_logic_vector(108 downto 0);
    iunit_exec_to_writeback_pipe_write_req : out  std_logic_vector(0 downto 0);
    iunit_exec_to_writeback_pipe_write_ack : in   std_logic_vector(0 downto 0);
    iunit_exec_to_writeback_pipe_write_data : out  std_logic_vector(125 downto 0);
    teu_iunit_to_stream_corrector_pipe_write_req : out  std_logic_vector(0 downto 0);
    teu_iunit_to_stream_corrector_pipe_write_ack : in   std_logic_vector(0 downto 0);
    teu_iunit_to_stream_corrector_pipe_write_data : out  std_logic_vector(89 downto 0);
    teu_iunit_trap_to_fpunit_pipe_write_req : out  std_logic_vector(0 downto 0);
    teu_iunit_trap_to_fpunit_pipe_write_ack : in   std_logic_vector(0 downto 0);
    teu_iunit_trap_to_fpunit_pipe_write_data : out  std_logic_vector(12 downto 0);
    teu_iunit_trap_to_loadstore_pipe_write_req : out  std_logic_vector(0 downto 0);
    teu_iunit_trap_to_loadstore_pipe_write_ack : in   std_logic_vector(0 downto 0);
    teu_iunit_trap_to_loadstore_pipe_write_data : out  std_logic_vector(0 downto 0);
    i32_div_call_reqs : out  std_logic_vector(0 downto 0);
    i32_div_call_acks : in   std_logic_vector(0 downto 0);
    i32_div_call_data : out  std_logic_vector(97 downto 0);
    i32_div_call_tag  :  out  std_logic_vector(0 downto 0);
    i32_div_return_reqs : out  std_logic_vector(0 downto 0);
    i32_div_return_acks : in   std_logic_vector(0 downto 0);
    i32_div_return_data : in   std_logic_vector(35 downto 0);
    i32_div_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity iu_exec_daemon;
architecture iu_exec_daemon_arch of iu_exec_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal iu_exec_daemon_CP_1081_start: Boolean;
  signal iu_exec_daemon_CP_1081_symbol: Boolean;
  -- volatile/operator module components. 
  component decode_alu_exec_control_word_Volatile is -- 
    port ( -- 
      cw : in  std_logic_vector(54 downto 0);
      cti : out  std_logic_vector(0 downto 0);
      is_call : out  std_logic_vector(0 downto 0);
      is_jmpl : out  std_logic_vector(0 downto 0);
      is_rett : out  std_logic_vector(0 downto 0);
      is_bicc : out  std_logic_vector(0 downto 0);
      is_fbfcc : out  std_logic_vector(0 downto 0);
      is_cbccc : out  std_logic_vector(0 downto 0);
      is_ticc : out  std_logic_vector(0 downto 0);
      annul_flag : out  std_logic_vector(0 downto 0);
      br_cond : out  std_logic_vector(3 downto 0);
      alu : out  std_logic_vector(0 downto 0);
      use_alu_add : out  std_logic_vector(0 downto 0);
      is_alu_sub : out  std_logic_vector(0 downto 0);
      is_alu_mul : out  std_logic_vector(0 downto 0);
      is_alu_mulscc : out  std_logic_vector(0 downto 0);
      is_alu_div : out  std_logic_vector(0 downto 0);
      is_alu_sll : out  std_logic_vector(0 downto 0);
      is_alu_srl : out  std_logic_vector(0 downto 0);
      is_alu_sra : out  std_logic_vector(0 downto 0);
      is_alu_and : out  std_logic_vector(0 downto 0);
      is_alu_or : out  std_logic_vector(0 downto 0);
      use_alu_xor : out  std_logic_vector(0 downto 0);
      is_alu_xnor : out  std_logic_vector(0 downto 0);
      signed_mul_div : out  std_logic_vector(0 downto 0);
      negate_second_operand : out  std_logic_vector(0 downto 0);
      with_carry : out  std_logic_vector(0 downto 0);
      set_cc : out  std_logic_vector(0 downto 0);
      tagged_alu_op : out  std_logic_vector(0 downto 0);
      trap_on_overflow : out  std_logic_vector(0 downto 0);
      misc : out  std_logic_vector(0 downto 0);
      is_sethi : out  std_logic_vector(0 downto 0);
      write_psr : out  std_logic_vector(0 downto 0);
      write_wim : out  std_logic_vector(0 downto 0);
      write_tbr : out  std_logic_vector(0 downto 0);
      write_y : out  std_logic_vector(0 downto 0);
      write_asr : out  std_logic_vector(0 downto 0);
      read_psr : out  std_logic_vector(0 downto 0);
      read_wim : out  std_logic_vector(0 downto 0);
      read_tbr : out  std_logic_vector(0 downto 0);
      read_y : out  std_logic_vector(0 downto 0);
      read_asr : out  std_logic_vector(0 downto 0);
      asr_id : out  std_logic_vector(4 downto 0);
      is_save : out  std_logic_vector(0 downto 0);
      is_restore : out  std_logic_vector(0 downto 0);
      dti : out  std_logic_vector(0 downto 0);
      is_iu_dti : out  std_logic_vector(0 downto 0);
      is_load_to_debug : out  std_logic_vector(0 downto 0);
      is_store_to_debug : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component i32_add_sub_Volatile is -- 
    port ( -- 
      subtract_flag : in  std_logic_vector(0 downto 0);
      with_carry : in  std_logic_vector(0 downto 0);
      set_cc : in  std_logic_vector(0 downto 0);
      tagged_op : in  std_logic_vector(0 downto 0);
      trap_on_ovflow : in  std_logic_vector(0 downto 0);
      Ni : in  std_logic_vector(0 downto 0);
      Zi : in  std_logic_vector(0 downto 0);
      Vi : in  std_logic_vector(0 downto 0);
      Ci : in  std_logic_vector(0 downto 0);
      x : in  std_logic_vector(31 downto 0);
      y : in  std_logic_vector(31 downto 0);
      result : out  std_logic_vector(31 downto 0);
      No : out  std_logic_vector(0 downto 0);
      Zo : out  std_logic_vector(0 downto 0);
      Vo : out  std_logic_vector(0 downto 0);
      Co : out  std_logic_vector(0 downto 0);
      overflow_trap : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component exec_cti_instruction_Volatile is -- 
    port ( -- 
      exec_call : in  std_logic_vector(0 downto 0);
      exec_rett : in  std_logic_vector(0 downto 0);
      exec_jmpl : in  std_logic_vector(0 downto 0);
      exec_ticc : in  std_logic_vector(0 downto 0);
      br_cond : in  std_logic_vector(3 downto 0);
      annul_flag : in  std_logic_vector(0 downto 0);
      pc : in  std_logic_vector(31 downto 0);
      alu_result : in  std_logic_vector(31 downto 0);
      psr : in  std_logic_vector(31 downto 0);
      wim : in  std_logic_vector(31 downto 0);
      cti_trap_status : out  std_logic_vector(0 downto 0);
      cti_ticc_trap_type : out  std_logic_vector(6 downto 0);
      cti_trap_instr_trap : out  std_logic_vector(0 downto 0);
      cti_illegal_instr_trap : out  std_logic_vector(0 downto 0);
      cti_privileged_instr_trap : out  std_logic_vector(0 downto 0);
      cti_window_underflow_trap : out  std_logic_vector(0 downto 0);
      cti_mem_address_not_aligned_trap : out  std_logic_vector(0 downto 0);
      cti_processor_error_mode : out  std_logic_vector(0 downto 0);
      cti_br_taken : out  std_logic_vector(0 downto 0);
      cti_next_psr : out  std_logic_vector(31 downto 0);
      cti_annul_next : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component i32_div is -- 
    generic (tag_length : integer); 
    port ( -- 
      signed_div : in  std_logic_vector(0 downto 0);
      set_cc : in  std_logic_vector(0 downto 0);
      y_in : in  std_logic_vector(31 downto 0);
      dividend : in  std_logic_vector(31 downto 0);
      divisor : in  std_logic_vector(31 downto 0);
      result : out  std_logic_vector(31 downto 0);
      No : out  std_logic_vector(0 downto 0);
      Zo : out  std_logic_vector(0 downto 0);
      Vo : out  std_logic_vector(0 downto 0);
      Co : out  std_logic_vector(0 downto 0);
      u64_true_divide_revised_call_reqs : out  std_logic_vector(0 downto 0);
      u64_true_divide_revised_call_acks : in   std_logic_vector(0 downto 0);
      u64_true_divide_revised_call_data : out  std_logic_vector(95 downto 0);
      u64_true_divide_revised_call_tag  :  out  std_logic_vector(0 downto 0);
      u64_true_divide_revised_return_reqs : out  std_logic_vector(0 downto 0);
      u64_true_divide_revised_return_acks : in   std_logic_vector(0 downto 0);
      u64_true_divide_revised_return_data : in   std_logic_vector(63 downto 0);
      u64_true_divide_revised_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component i32_mulscc_Volatile is -- 
    port ( -- 
      y_in : in  std_logic_vector(31 downto 0);
      A : in  std_logic_vector(31 downto 0);
      B : in  std_logic_vector(31 downto 0);
      Ni : in  std_logic_vector(0 downto 0);
      Zi : in  std_logic_vector(0 downto 0);
      Vi : in  std_logic_vector(0 downto 0);
      Ci : in  std_logic_vector(0 downto 0);
      y_out : out  std_logic_vector(31 downto 0);
      result : out  std_logic_vector(31 downto 0);
      No : out  std_logic_vector(0 downto 0);
      Zo : out  std_logic_vector(0 downto 0);
      Vo : out  std_logic_vector(0 downto 0);
      Co : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component restore_window_trap_Volatile is -- 
    port ( -- 
      psr : in  std_logic_vector(31 downto 0);
      wim : in  std_logic_vector(31 downto 0);
      uflow_trap : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- function library module [iu_umul32] component not printed.
  component i32_mul_calculate_sign_correction_Volatile is -- 
    port ( -- 
      signed_mul : in  std_logic_vector(0 downto 0);
      A : in  std_logic_vector(31 downto 0);
      B : in  std_logic_vector(31 downto 0);
      sign_correction : out  std_logic_vector(31 downto 0)-- 
    );
    -- 
  end component; 
  component i32_shift_Volatile is -- 
    port ( -- 
      is_sll : in  std_logic_vector(0 downto 0);
      is_srl : in  std_logic_vector(0 downto 0);
      is_sra : in  std_logic_vector(0 downto 0);
      x : in  std_logic_vector(31 downto 0);
      shift_amount : in  std_logic_vector(31 downto 0);
      result : out  std_logic_vector(31 downto 0)-- 
    );
    -- 
  end component; 
  component save_window_trap_Volatile is -- 
    port ( -- 
      psr : in  std_logic_vector(31 downto 0);
      wim : in  std_logic_vector(31 downto 0);
      ovflow_trap : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_inst_req_1 : boolean;
  signal W_exec_info_d_8377_inst_req_0 : boolean;
  signal do_while_stmt_8361_branch_req_0 : boolean;
  signal WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_inst_req_0 : boolean;
  signal W_exec_info_d_8377_inst_ack_0 : boolean;
  signal RPIPE_iunit_register_file_read_access_response_8375_inst_ack_1 : boolean;
  signal W_issue_mul_9416_delayed_1_0_9244_inst_ack_0 : boolean;
  signal WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_inst_req_1 : boolean;
  signal WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_inst_ack_1 : boolean;
  signal WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_inst_req_1 : boolean;
  signal W_issue_mul_9416_delayed_1_0_9244_inst_req_0 : boolean;
  signal CONCAT_u2_u4_9254_inst_req_0 : boolean;
  signal W_issue_mul_9416_delayed_1_0_9244_inst_ack_1 : boolean;
  signal WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_inst_ack_1 : boolean;
  signal WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_inst_req_0 : boolean;
  signal WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_inst_ack_1 : boolean;
  signal WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_inst_ack_0 : boolean;
  signal call_stmt_9223_call_req_1 : boolean;
  signal WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_inst_ack_0 : boolean;
  signal RPIPE_iunit_register_file_read_access_response_8375_inst_req_1 : boolean;
  signal CONCAT_u2_u4_9254_inst_req_1 : boolean;
  signal W_exec_info_d_8377_inst_req_1 : boolean;
  signal W_exec_info_d_8377_inst_ack_1 : boolean;
  signal WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_inst_req_1 : boolean;
  signal RPIPE_iunit_register_file_read_access_response_8375_inst_req_0 : boolean;
  signal WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_inst_ack_1 : boolean;
  signal W_issue_mul_9416_delayed_1_0_9244_inst_req_1 : boolean;
  signal CONCAT_u2_u4_9254_inst_ack_0 : boolean;
  signal RPIPE_iunit_register_file_read_access_response_8375_inst_ack_0 : boolean;
  signal call_stmt_9223_call_ack_0 : boolean;
  signal call_stmt_9223_call_req_0 : boolean;
  signal W_get_from_rfile_8647_delayed_1_0_8476_inst_ack_1 : boolean;
  signal W_issue_div_9432_delayed_1_0_9268_inst_ack_0 : boolean;
  signal RPIPE_teu_idispatch_to_iunit_exec_8364_inst_ack_1 : boolean;
  signal MUX_9296_inst_req_1 : boolean;
  signal MUX_9296_inst_ack_1 : boolean;
  signal W_get_from_rfile_8647_delayed_1_0_8476_inst_req_1 : boolean;
  signal W_issue_div_9432_delayed_1_0_9268_inst_req_0 : boolean;
  signal RPIPE_teu_idispatch_to_iunit_exec_8364_inst_req_1 : boolean;
  signal MUX_9296_inst_ack_0 : boolean;
  signal MUX_9296_inst_req_0 : boolean;
  signal W_issue_add_sub_9424_delayed_1_0_9256_inst_ack_1 : boolean;
  signal W_get_from_rfile_8647_delayed_1_0_8476_inst_ack_0 : boolean;
  signal WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_inst_ack_0 : boolean;
  signal CONCAT_u2_u4_9266_inst_ack_0 : boolean;
  signal CONCAT_u2_u4_9266_inst_req_0 : boolean;
  signal W_issue_add_sub_9424_delayed_1_0_9256_inst_ack_0 : boolean;
  signal W_issue_add_sub_9424_delayed_1_0_9256_inst_req_1 : boolean;
  signal W_issue_add_sub_9424_delayed_1_0_9256_inst_req_0 : boolean;
  signal RPIPE_teu_idispatch_to_iunit_exec_8364_inst_ack_0 : boolean;
  signal WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_inst_ack_0 : boolean;
  signal RPIPE_teu_idispatch_to_iunit_exec_8364_inst_req_0 : boolean;
  signal WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_inst_req_0 : boolean;
  signal W_get_from_rfile_8647_delayed_1_0_8476_inst_req_0 : boolean;
  signal WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_inst_req_0 : boolean;
  signal CONCAT_u2_u4_9266_inst_req_1 : boolean;
  signal CONCAT_u2_u4_9266_inst_ack_1 : boolean;
  signal CONCAT_u2_u4_9254_inst_ack_1 : boolean;
  signal call_stmt_9223_call_ack_1 : boolean;
  signal W_issue_div_9432_delayed_1_0_9268_inst_req_1 : boolean;
  signal W_issue_div_9432_delayed_1_0_9268_inst_ack_1 : boolean;
  signal slice_9318_inst_req_0 : boolean;
  signal slice_9318_inst_ack_0 : boolean;
  signal slice_9318_inst_req_1 : boolean;
  signal slice_9318_inst_ack_1 : boolean;
  signal slice_9322_inst_req_0 : boolean;
  signal slice_9322_inst_ack_0 : boolean;
  signal slice_9322_inst_req_1 : boolean;
  signal slice_9322_inst_ack_1 : boolean;
  signal W_issue_mul_9479_delayed_1_0_9331_inst_req_0 : boolean;
  signal W_issue_mul_9479_delayed_1_0_9331_inst_ack_0 : boolean;
  signal W_issue_mul_9479_delayed_1_0_9331_inst_req_1 : boolean;
  signal W_issue_mul_9479_delayed_1_0_9331_inst_ack_1 : boolean;
  signal W_i32_mul_result_9480_delayed_1_0_9334_inst_req_0 : boolean;
  signal W_i32_mul_result_9480_delayed_1_0_9334_inst_ack_0 : boolean;
  signal W_i32_mul_result_9480_delayed_1_0_9334_inst_req_1 : boolean;
  signal W_i32_mul_result_9480_delayed_1_0_9334_inst_ack_1 : boolean;
  signal MUX_9347_inst_req_0 : boolean;
  signal MUX_9347_inst_ack_0 : boolean;
  signal MUX_9347_inst_req_1 : boolean;
  signal MUX_9347_inst_ack_1 : boolean;
  signal W_issue_div_9491_delayed_1_0_9349_inst_req_0 : boolean;
  signal W_issue_div_9491_delayed_1_0_9349_inst_ack_0 : boolean;
  signal W_issue_div_9491_delayed_1_0_9349_inst_req_1 : boolean;
  signal W_issue_div_9491_delayed_1_0_9349_inst_ack_1 : boolean;
  signal OR_u32_u32_9361_inst_req_0 : boolean;
  signal OR_u32_u32_9361_inst_ack_0 : boolean;
  signal OR_u32_u32_9361_inst_req_1 : boolean;
  signal OR_u32_u32_9361_inst_ack_1 : boolean;
  signal OR_u32_u32_9382_inst_req_0 : boolean;
  signal OR_u32_u32_9382_inst_ack_0 : boolean;
  signal OR_u32_u32_9382_inst_req_1 : boolean;
  signal OR_u32_u32_9382_inst_ack_1 : boolean;
  signal OR_u1_u1_9437_inst_req_0 : boolean;
  signal OR_u1_u1_9437_inst_ack_0 : boolean;
  signal OR_u1_u1_9437_inst_req_1 : boolean;
  signal OR_u1_u1_9437_inst_ack_1 : boolean;
  signal W_psr_9567_delayed_1_0_9439_inst_req_0 : boolean;
  signal W_psr_9567_delayed_1_0_9439_inst_ack_0 : boolean;
  signal W_psr_9567_delayed_1_0_9439_inst_req_1 : boolean;
  signal W_psr_9567_delayed_1_0_9439_inst_ack_1 : boolean;
  signal W_exec_rett_9568_delayed_1_0_9442_inst_req_0 : boolean;
  signal W_exec_rett_9568_delayed_1_0_9442_inst_ack_0 : boolean;
  signal W_exec_rett_9568_delayed_1_0_9442_inst_req_1 : boolean;
  signal W_exec_rett_9568_delayed_1_0_9442_inst_ack_1 : boolean;
  signal W_cti_next_psr_9569_delayed_1_0_9445_inst_req_0 : boolean;
  signal W_cti_next_psr_9569_delayed_1_0_9445_inst_ack_0 : boolean;
  signal W_cti_next_psr_9569_delayed_1_0_9445_inst_req_1 : boolean;
  signal W_cti_next_psr_9569_delayed_1_0_9445_inst_ack_1 : boolean;
  signal W_write_psr_9570_delayed_1_0_9448_inst_req_0 : boolean;
  signal W_write_psr_9570_delayed_1_0_9448_inst_ack_0 : boolean;
  signal W_write_psr_9570_delayed_1_0_9448_inst_req_1 : boolean;
  signal W_write_psr_9570_delayed_1_0_9448_inst_ack_1 : boolean;
  signal W_i32_xor_result_9571_delayed_1_0_9451_inst_req_0 : boolean;
  signal W_i32_xor_result_9571_delayed_1_0_9451_inst_ack_0 : boolean;
  signal W_i32_xor_result_9571_delayed_1_0_9451_inst_req_1 : boolean;
  signal W_i32_xor_result_9571_delayed_1_0_9451_inst_ack_1 : boolean;
  signal OR_u1_u1_9465_inst_req_0 : boolean;
  signal OR_u1_u1_9465_inst_ack_0 : boolean;
  signal OR_u1_u1_9465_inst_req_1 : boolean;
  signal OR_u1_u1_9465_inst_ack_1 : boolean;
  signal W_psr_9584_delayed_1_0_9467_inst_req_0 : boolean;
  signal W_psr_9584_delayed_1_0_9467_inst_ack_0 : boolean;
  signal W_psr_9584_delayed_1_0_9467_inst_req_1 : boolean;
  signal W_psr_9584_delayed_1_0_9467_inst_ack_1 : boolean;
  signal WPIPE_teu_iunit_to_stream_corrector_9734_inst_req_0 : boolean;
  signal WPIPE_teu_iunit_to_stream_corrector_9734_inst_ack_0 : boolean;
  signal WPIPE_teu_iunit_to_stream_corrector_9734_inst_req_1 : boolean;
  signal WPIPE_teu_iunit_to_stream_corrector_9734_inst_ack_1 : boolean;
  signal CONCAT_u12_u14_9763_inst_req_0 : boolean;
  signal CONCAT_u12_u14_9763_inst_ack_0 : boolean;
  signal CONCAT_u12_u14_9763_inst_req_1 : boolean;
  signal CONCAT_u12_u14_9763_inst_ack_1 : boolean;
  signal CONCAT_u15_u16_9768_inst_req_0 : boolean;
  signal CONCAT_u15_u16_9768_inst_ack_0 : boolean;
  signal CONCAT_u15_u16_9768_inst_req_1 : boolean;
  signal CONCAT_u15_u16_9768_inst_ack_1 : boolean;
  signal W_updated_y_9874_delayed_1_0_9770_inst_req_0 : boolean;
  signal W_updated_y_9874_delayed_1_0_9770_inst_ack_0 : boolean;
  signal W_updated_y_9874_delayed_1_0_9770_inst_req_1 : boolean;
  signal W_updated_y_9874_delayed_1_0_9770_inst_ack_1 : boolean;
  signal W_send_to_wb_9880_delayed_1_0_9784_inst_req_0 : boolean;
  signal W_send_to_wb_9880_delayed_1_0_9784_inst_ack_0 : boolean;
  signal W_send_to_wb_9880_delayed_1_0_9784_inst_req_1 : boolean;
  signal W_send_to_wb_9880_delayed_1_0_9784_inst_ack_1 : boolean;
  signal WPIPE_iunit_exec_to_writeback_9788_inst_req_0 : boolean;
  signal WPIPE_iunit_exec_to_writeback_9788_inst_ack_0 : boolean;
  signal WPIPE_iunit_exec_to_writeback_9788_inst_req_1 : boolean;
  signal WPIPE_iunit_exec_to_writeback_9788_inst_ack_1 : boolean;
  signal WPIPE_teu_iunit_trap_to_loadstore_9821_inst_req_0 : boolean;
  signal WPIPE_teu_iunit_trap_to_loadstore_9821_inst_ack_0 : boolean;
  signal WPIPE_teu_iunit_trap_to_loadstore_9821_inst_req_1 : boolean;
  signal WPIPE_teu_iunit_trap_to_loadstore_9821_inst_ack_1 : boolean;
  signal WPIPE_teu_iunit_trap_to_fpunit_9840_inst_req_0 : boolean;
  signal WPIPE_teu_iunit_trap_to_fpunit_9840_inst_ack_0 : boolean;
  signal WPIPE_teu_iunit_trap_to_fpunit_9840_inst_req_1 : boolean;
  signal WPIPE_teu_iunit_trap_to_fpunit_9840_inst_ack_1 : boolean;
  signal do_while_stmt_8361_branch_ack_0 : boolean;
  signal do_while_stmt_8361_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "iu_exec_daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  iu_exec_daemon_CP_1081_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "iu_exec_daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= iu_exec_daemon_CP_1081_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= iu_exec_daemon_CP_1081_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= iu_exec_daemon_CP_1081_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  iu_exec_daemon_CP_1081: Block -- control-path 
    signal iu_exec_daemon_CP_1081_elements: BooleanArray(154 downto 0);
    -- 
  begin -- 
    iu_exec_daemon_CP_1081_elements(0) <= iu_exec_daemon_CP_1081_start;
    iu_exec_daemon_CP_1081_symbol <= iu_exec_daemon_CP_1081_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_8360/branch_block_stmt_8360__entry__
      -- CP-element group 0: 	 branch_block_stmt_8360/do_while_stmt_8361__entry__
      -- CP-element group 0: 	 branch_block_stmt_8360/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	154 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_8360/do_while_stmt_8361__exit__
      -- CP-element group 1: 	 branch_block_stmt_8360/$exit
      -- CP-element group 1: 	 branch_block_stmt_8360/branch_block_stmt_8360__exit__
      -- CP-element group 1: 	 $exit
      -- 
    iu_exec_daemon_CP_1081_elements(1) <= iu_exec_daemon_CP_1081_elements(154);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_8360/do_while_stmt_8361/$entry
      -- CP-element group 2: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361__entry__
      -- 
    iu_exec_daemon_CP_1081_elements(2) <= iu_exec_daemon_CP_1081_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	154 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361__exit__
      -- 
    -- Element group iu_exec_daemon_CP_1081_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_8360/do_while_stmt_8361/loop_back
      -- 
    -- Element group iu_exec_daemon_CP_1081_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	150 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	152 
    -- CP-element group 5: 	153 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_8360/do_while_stmt_8361/condition_done
      -- CP-element group 5: 	 branch_block_stmt_8360/do_while_stmt_8361/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_8360/do_while_stmt_8361/loop_taken/$entry
      -- 
    iu_exec_daemon_CP_1081_elements(5) <= iu_exec_daemon_CP_1081_elements(150);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	151 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_8360/do_while_stmt_8361/loop_body_done
      -- 
    iu_exec_daemon_CP_1081_elements(6) <= iu_exec_daemon_CP_1081_elements(151);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/back_edge_to_loop_body
      -- 
    iu_exec_daemon_CP_1081_elements(7) <= iu_exec_daemon_CP_1081_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/first_time_through_loop_body
      -- 
    iu_exec_daemon_CP_1081_elements(8) <= iu_exec_daemon_CP_1081_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	150 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/loop_body_start
      -- 
    -- Element group iu_exec_daemon_CP_1081_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_teu_idispatch_to_iunit_exec_8364_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_teu_idispatch_to_iunit_exec_8364_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_teu_idispatch_to_iunit_exec_8364_Sample/$entry
      -- 
    rr_1114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(10), ack => RPIPE_teu_idispatch_to_iunit_exec_8364_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(9) & iu_exec_daemon_CP_1081_elements(13);
      gj_iu_exec_daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	19 
    -- CP-element group 11: 	22 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_teu_idispatch_to_iunit_exec_8364_update_start_
      -- CP-element group 11: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_teu_idispatch_to_iunit_exec_8364_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_teu_idispatch_to_iunit_exec_8364_Update/$entry
      -- 
    cr_1119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(11), ack => RPIPE_teu_idispatch_to_iunit_exec_8364_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(12) & iu_exec_daemon_CP_1081_elements(16) & iu_exec_daemon_CP_1081_elements(19) & iu_exec_daemon_CP_1081_elements(22);
      gj_iu_exec_daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_teu_idispatch_to_iunit_exec_8364_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_teu_idispatch_to_iunit_exec_8364_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_teu_idispatch_to_iunit_exec_8364_Sample/$exit
      -- 
    ra_1115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_teu_idispatch_to_iunit_exec_8364_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	22 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8379_Sample/req
      -- CP-element group 13: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8478_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8379_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8478_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_teu_idispatch_to_iunit_exec_8364_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_teu_idispatch_to_iunit_exec_8364_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8478_Sample/req
      -- CP-element group 13: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8379_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_teu_idispatch_to_iunit_exec_8364_update_completed_
      -- 
    ca_1120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_teu_idispatch_to_iunit_exec_8364_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(13)); -- 
    req_1142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(13), ack => W_exec_info_d_8377_inst_req_0); -- 
    req_1156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(13), ack => W_get_from_rfile_8647_delayed_1_0_8476_inst_req_0); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_iunit_register_file_read_access_response_8375_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_iunit_register_file_read_access_response_8375_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_iunit_register_file_read_access_response_8375_sample_start_
      -- 
    rr_1128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(14), ack => RPIPE_iunit_register_file_read_access_response_8375_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(13) & iu_exec_daemon_CP_1081_elements(17);
      gj_iu_exec_daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	95 
    -- CP-element group 15: 	68 
    -- CP-element group 15: 	91 
    -- CP-element group 15: 	79 
    -- CP-element group 15: 	87 
    -- CP-element group 15: 	83 
    -- CP-element group 15: 	121 
    -- CP-element group 15: 	124 
    -- CP-element group 15: 	128 
    -- CP-element group 15: 	132 
    -- CP-element group 15: 	136 
    -- CP-element group 15: 	145 
    -- CP-element group 15: 	148 
    -- CP-element group 15: 	75 
    -- CP-element group 15: 	113 
    -- CP-element group 15: 	117 
    -- CP-element group 15: 	106 
    -- CP-element group 15: 	99 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	31 
    -- CP-element group 15: 	34 
    -- CP-element group 15: 	38 
    -- CP-element group 15: 	45 
    -- CP-element group 15: 	52 
    -- CP-element group 15: 	56 
    -- CP-element group 15: 	60 
    -- CP-element group 15: 	64 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_iunit_register_file_read_access_response_8375_update_start_
      -- CP-element group 15: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_iunit_register_file_read_access_response_8375_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_iunit_register_file_read_access_response_8375_Update/cr
      -- 
    cr_1133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(15), ack => RPIPE_iunit_register_file_read_access_response_8375_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 28) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1);
      constant place_markings: IntegerArray(0 to 28)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1);
      constant place_delays: IntegerArray(0 to 28) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 29); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(16) & iu_exec_daemon_CP_1081_elements(95) & iu_exec_daemon_CP_1081_elements(68) & iu_exec_daemon_CP_1081_elements(91) & iu_exec_daemon_CP_1081_elements(79) & iu_exec_daemon_CP_1081_elements(87) & iu_exec_daemon_CP_1081_elements(83) & iu_exec_daemon_CP_1081_elements(121) & iu_exec_daemon_CP_1081_elements(124) & iu_exec_daemon_CP_1081_elements(128) & iu_exec_daemon_CP_1081_elements(132) & iu_exec_daemon_CP_1081_elements(136) & iu_exec_daemon_CP_1081_elements(145) & iu_exec_daemon_CP_1081_elements(148) & iu_exec_daemon_CP_1081_elements(75) & iu_exec_daemon_CP_1081_elements(113) & iu_exec_daemon_CP_1081_elements(117) & iu_exec_daemon_CP_1081_elements(106) & iu_exec_daemon_CP_1081_elements(99) & iu_exec_daemon_CP_1081_elements(25) & iu_exec_daemon_CP_1081_elements(28) & iu_exec_daemon_CP_1081_elements(31) & iu_exec_daemon_CP_1081_elements(34) & iu_exec_daemon_CP_1081_elements(38) & iu_exec_daemon_CP_1081_elements(45) & iu_exec_daemon_CP_1081_elements(52) & iu_exec_daemon_CP_1081_elements(56) & iu_exec_daemon_CP_1081_elements(60) & iu_exec_daemon_CP_1081_elements(64);
      gj_iu_exec_daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 29, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_iunit_register_file_read_access_response_8375_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_iunit_register_file_read_access_response_8375_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_iunit_register_file_read_access_response_8375_sample_completed_
      -- 
    ra_1129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_iunit_register_file_read_access_response_8375_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	97 
    -- CP-element group 17: 	73 
    -- CP-element group 17: 	81 
    -- CP-element group 17: 	85 
    -- CP-element group 17: 	89 
    -- CP-element group 17: 	93 
    -- CP-element group 17: 	77 
    -- CP-element group 17: 	119 
    -- CP-element group 17: 	123 
    -- CP-element group 17: 	126 
    -- CP-element group 17: 	130 
    -- CP-element group 17: 	134 
    -- CP-element group 17: 	144 
    -- CP-element group 17: 	147 
    -- CP-element group 17: 	111 
    -- CP-element group 17: 	115 
    -- CP-element group 17: 	104 
    -- CP-element group 17: 	24 
    -- CP-element group 17: 	27 
    -- CP-element group 17: 	30 
    -- CP-element group 17: 	33 
    -- CP-element group 17: 	36 
    -- CP-element group 17: 	43 
    -- CP-element group 17: 	50 
    -- CP-element group 17: 	54 
    -- CP-element group 17: 	58 
    -- CP-element group 17: 	62 
    -- CP-element group 17: 	66 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_iunit_register_file_read_access_response_8375_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_iunit_register_file_read_access_response_8375_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/RPIPE_iunit_register_file_read_access_response_8375_Update/ca
      -- 
    ca_1134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_iunit_register_file_read_access_response_8375_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	95 
    -- CP-element group 18: 	71 
    -- CP-element group 18: 	91 
    -- CP-element group 18: 	79 
    -- CP-element group 18: 	87 
    -- CP-element group 18: 	83 
    -- CP-element group 18: 	124 
    -- CP-element group 18: 	128 
    -- CP-element group 18: 	132 
    -- CP-element group 18: 	136 
    -- CP-element group 18: 	139 
    -- CP-element group 18: 	145 
    -- CP-element group 18: 	148 
    -- CP-element group 18: 	75 
    -- CP-element group 18: 	113 
    -- CP-element group 18: 	117 
    -- CP-element group 18: 	106 
    -- CP-element group 18: 	109 
    -- CP-element group 18: 	102 
    -- CP-element group 18: 	28 
    -- CP-element group 18: 	31 
    -- CP-element group 18: 	34 
    -- CP-element group 18: 	38 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	45 
    -- CP-element group 18: 	48 
    -- CP-element group 18: 	52 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	60 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8379_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8379_update_start_
      -- CP-element group 18: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8379_Update/req
      -- 
    req_1147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(18), ack => W_exec_info_d_8377_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 28) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1);
      constant place_markings: IntegerArray(0 to 28)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1);
      constant place_delays: IntegerArray(0 to 28) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 29); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(95) & iu_exec_daemon_CP_1081_elements(71) & iu_exec_daemon_CP_1081_elements(91) & iu_exec_daemon_CP_1081_elements(79) & iu_exec_daemon_CP_1081_elements(87) & iu_exec_daemon_CP_1081_elements(83) & iu_exec_daemon_CP_1081_elements(124) & iu_exec_daemon_CP_1081_elements(128) & iu_exec_daemon_CP_1081_elements(132) & iu_exec_daemon_CP_1081_elements(136) & iu_exec_daemon_CP_1081_elements(139) & iu_exec_daemon_CP_1081_elements(145) & iu_exec_daemon_CP_1081_elements(148) & iu_exec_daemon_CP_1081_elements(75) & iu_exec_daemon_CP_1081_elements(113) & iu_exec_daemon_CP_1081_elements(117) & iu_exec_daemon_CP_1081_elements(106) & iu_exec_daemon_CP_1081_elements(109) & iu_exec_daemon_CP_1081_elements(102) & iu_exec_daemon_CP_1081_elements(28) & iu_exec_daemon_CP_1081_elements(31) & iu_exec_daemon_CP_1081_elements(34) & iu_exec_daemon_CP_1081_elements(38) & iu_exec_daemon_CP_1081_elements(41) & iu_exec_daemon_CP_1081_elements(45) & iu_exec_daemon_CP_1081_elements(48) & iu_exec_daemon_CP_1081_elements(52) & iu_exec_daemon_CP_1081_elements(56) & iu_exec_daemon_CP_1081_elements(60);
      gj_iu_exec_daemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 29, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	11 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8379_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8379_Sample/ack
      -- CP-element group 19: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8379_Sample/$exit
      -- 
    ack_1143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_exec_info_d_8377_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	71 
    -- CP-element group 20: 	73 
    -- CP-element group 20: 	81 
    -- CP-element group 20: 	85 
    -- CP-element group 20: 	89 
    -- CP-element group 20: 	93 
    -- CP-element group 20: 	77 
    -- CP-element group 20: 	123 
    -- CP-element group 20: 	126 
    -- CP-element group 20: 	130 
    -- CP-element group 20: 	134 
    -- CP-element group 20: 	139 
    -- CP-element group 20: 	144 
    -- CP-element group 20: 	147 
    -- CP-element group 20: 	111 
    -- CP-element group 20: 	115 
    -- CP-element group 20: 	104 
    -- CP-element group 20: 	109 
    -- CP-element group 20: 	102 
    -- CP-element group 20: 	27 
    -- CP-element group 20: 	30 
    -- CP-element group 20: 	33 
    -- CP-element group 20: 	36 
    -- CP-element group 20: 	41 
    -- CP-element group 20: 	43 
    -- CP-element group 20: 	48 
    -- CP-element group 20: 	50 
    -- CP-element group 20: 	54 
    -- CP-element group 20: 	58 
    -- CP-element group 20:  members (21) 
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8379_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9246_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9246_Sample/req
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9258_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8379_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8379_Update/ack
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9246_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9258_Sample/req
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9258_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9333_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9333_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9333_Sample/req
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9444_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9444_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9444_Sample/req
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9450_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9450_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9450_Sample/req
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9786_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9786_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9786_Sample/req
      -- 
    ack_1148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_exec_info_d_8377_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(20)); -- 
    req_1352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(20), ack => W_issue_mul_9479_delayed_1_0_9331_inst_req_0); -- 
    req_1604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(20), ack => W_send_to_wb_9880_delayed_1_0_9784_inst_req_0); -- 
    req_1492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(20), ack => W_write_psr_9570_delayed_1_0_9448_inst_req_0); -- 
    req_1464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(20), ack => W_exec_rett_9568_delayed_1_0_9442_inst_req_0); -- 
    req_1240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(20), ack => W_issue_mul_9416_delayed_1_0_9244_inst_req_0); -- 
    req_1268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(20), ack => W_issue_add_sub_9424_delayed_1_0_9256_inst_req_0); -- 
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	95 
    -- CP-element group 21: 	68 
    -- CP-element group 21: 	91 
    -- CP-element group 21: 	79 
    -- CP-element group 21: 	87 
    -- CP-element group 21: 	83 
    -- CP-element group 21: 	121 
    -- CP-element group 21: 	124 
    -- CP-element group 21: 	128 
    -- CP-element group 21: 	132 
    -- CP-element group 21: 	136 
    -- CP-element group 21: 	145 
    -- CP-element group 21: 	148 
    -- CP-element group 21: 	75 
    -- CP-element group 21: 	113 
    -- CP-element group 21: 	117 
    -- CP-element group 21: 	106 
    -- CP-element group 21: 	99 
    -- CP-element group 21: 	25 
    -- CP-element group 21: 	28 
    -- CP-element group 21: 	31 
    -- CP-element group 21: 	34 
    -- CP-element group 21: 	38 
    -- CP-element group 21: 	45 
    -- CP-element group 21: 	52 
    -- CP-element group 21: 	56 
    -- CP-element group 21: 	60 
    -- CP-element group 21: 	64 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8478_update_start_
      -- CP-element group 21: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8478_Update/req
      -- CP-element group 21: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8478_Update/$entry
      -- 
    req_1161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(21), ack => W_get_from_rfile_8647_delayed_1_0_8476_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 27) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1);
      constant place_markings: IntegerArray(0 to 27)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1);
      constant place_delays: IntegerArray(0 to 27) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 28); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(95) & iu_exec_daemon_CP_1081_elements(68) & iu_exec_daemon_CP_1081_elements(91) & iu_exec_daemon_CP_1081_elements(79) & iu_exec_daemon_CP_1081_elements(87) & iu_exec_daemon_CP_1081_elements(83) & iu_exec_daemon_CP_1081_elements(121) & iu_exec_daemon_CP_1081_elements(124) & iu_exec_daemon_CP_1081_elements(128) & iu_exec_daemon_CP_1081_elements(132) & iu_exec_daemon_CP_1081_elements(136) & iu_exec_daemon_CP_1081_elements(145) & iu_exec_daemon_CP_1081_elements(148) & iu_exec_daemon_CP_1081_elements(75) & iu_exec_daemon_CP_1081_elements(113) & iu_exec_daemon_CP_1081_elements(117) & iu_exec_daemon_CP_1081_elements(106) & iu_exec_daemon_CP_1081_elements(99) & iu_exec_daemon_CP_1081_elements(25) & iu_exec_daemon_CP_1081_elements(28) & iu_exec_daemon_CP_1081_elements(31) & iu_exec_daemon_CP_1081_elements(34) & iu_exec_daemon_CP_1081_elements(38) & iu_exec_daemon_CP_1081_elements(45) & iu_exec_daemon_CP_1081_elements(52) & iu_exec_daemon_CP_1081_elements(56) & iu_exec_daemon_CP_1081_elements(60) & iu_exec_daemon_CP_1081_elements(64);
      gj_iu_exec_daemon_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 28, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	13 
    -- CP-element group 22: successors 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	11 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8478_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8478_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8478_Sample/ack
      -- 
    ack_1157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_get_from_rfile_8647_delayed_1_0_8476_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	97 
    -- CP-element group 23: 	73 
    -- CP-element group 23: 	81 
    -- CP-element group 23: 	85 
    -- CP-element group 23: 	89 
    -- CP-element group 23: 	93 
    -- CP-element group 23: 	77 
    -- CP-element group 23: 	119 
    -- CP-element group 23: 	123 
    -- CP-element group 23: 	126 
    -- CP-element group 23: 	130 
    -- CP-element group 23: 	134 
    -- CP-element group 23: 	144 
    -- CP-element group 23: 	147 
    -- CP-element group 23: 	111 
    -- CP-element group 23: 	115 
    -- CP-element group 23: 	104 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	27 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	33 
    -- CP-element group 23: 	36 
    -- CP-element group 23: 	43 
    -- CP-element group 23: 	50 
    -- CP-element group 23: 	54 
    -- CP-element group 23: 	58 
    -- CP-element group 23: 	62 
    -- CP-element group 23: 	66 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8478_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8478_Update/ack
      -- CP-element group 23: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_8478_Update/$exit
      -- 
    ack_1162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_get_from_rfile_8647_delayed_1_0_8476_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	17 
    -- CP-element group 24: 	23 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_Sample/req
      -- 
    req_1170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(24), ack => WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(23) & iu_exec_daemon_CP_1081_elements(26);
      gj_iu_exec_daemon_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: 	21 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_update_start_
      -- CP-element group 25: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_Sample/ack
      -- CP-element group 25: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_Update/req
      -- 
    ack_1171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(25)); -- 
    req_1175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(25), ack => WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	151 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_Update/ack
      -- 
    ack_1176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	17 
    -- CP-element group 27: 	20 
    -- CP-element group 27: 	23 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_Sample/req
      -- CP-element group 27: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_Sample/$entry
      -- 
    req_1184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(27), ack => WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23) & iu_exec_daemon_CP_1081_elements(29);
      gj_iu_exec_daemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: 	18 
    -- CP-element group 28: 	21 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_Update/req
      -- CP-element group 28: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_update_start_
      -- CP-element group 28: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_Sample/$exit
      -- 
    ack_1185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(28)); -- 
    req_1189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(28), ack => WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_inst_req_1); -- 
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	151 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_Update/ack
      -- CP-element group 29: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_update_completed_
      -- 
    ack_1190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: 	20 
    -- CP-element group 30: 	23 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_Sample/req
      -- CP-element group 30: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_Sample/$entry
      -- 
    req_1198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(30), ack => WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23) & iu_exec_daemon_CP_1081_elements(32);
      gj_iu_exec_daemon_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	15 
    -- CP-element group 31: 	18 
    -- CP-element group 31: 	21 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_Update/req
      -- CP-element group 31: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_update_start_
      -- CP-element group 31: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_Sample/ack
      -- CP-element group 31: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_Sample/$exit
      -- 
    ack_1199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(31)); -- 
    req_1203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(31), ack => WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_inst_req_1); -- 
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	151 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_Update/ack
      -- 
    ack_1204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	17 
    -- CP-element group 33: 	20 
    -- CP-element group 33: 	23 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_Sample/req
      -- CP-element group 33: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_sample_start_
      -- 
    req_1212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(33), ack => WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23) & iu_exec_daemon_CP_1081_elements(35);
      gj_iu_exec_daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	15 
    -- CP-element group 34: 	18 
    -- CP-element group 34: 	21 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_Update/req
      -- CP-element group 34: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_Sample/ack
      -- CP-element group 34: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_update_start_
      -- CP-element group 34: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_Update/$entry
      -- 
    ack_1213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(34)); -- 
    req_1217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(34), ack => WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	151 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_Update/ack
      -- CP-element group 35: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_Update/$exit
      -- 
    ack_1218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	17 
    -- CP-element group 36: 	20 
    -- CP-element group 36: 	23 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/call_stmt_9223_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/call_stmt_9223_Sample/crr
      -- CP-element group 36: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/call_stmt_9223_Sample/$entry
      -- 
    crr_1226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(36), ack => call_stmt_9223_call_req_0); -- 
    iu_exec_daemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	142 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/call_stmt_9223_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/call_stmt_9223_Update/ccr
      -- CP-element group 37: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/call_stmt_9223_update_start_
      -- 
    ccr_1231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(37), ack => call_stmt_9223_call_req_1); -- 
    iu_exec_daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	15 
    -- CP-element group 38: 	18 
    -- CP-element group 38: 	21 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/call_stmt_9223_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/call_stmt_9223_Sample/cra
      -- CP-element group 38: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/call_stmt_9223_Sample/$exit
      -- 
    cra_1227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_9223_call_ack_0, ack => iu_exec_daemon_CP_1081_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	141 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/call_stmt_9223_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/call_stmt_9223_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/call_stmt_9223_Update/cca
      -- 
    cca_1232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_9223_call_ack_1, ack => iu_exec_daemon_CP_1081_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	142 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9246_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9246_update_start_
      -- CP-element group 40: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9246_Update/req
      -- 
    req_1245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(40), ack => W_issue_mul_9416_delayed_1_0_9244_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	20 
    -- CP-element group 41: successors 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	18 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9246_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9246_Sample/ack
      -- CP-element group 41: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9246_sample_completed_
      -- 
    ack_1241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_issue_mul_9416_delayed_1_0_9244_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	141 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9246_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9246_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9246_update_completed_
      -- 
    ack_1246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_issue_mul_9416_delayed_1_0_9244_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(42)); -- 
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	17 
    -- CP-element group 43: 	20 
    -- CP-element group 43: 	23 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9254_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9254_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9254_sample_start_
      -- 
    rr_1254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(43), ack => CONCAT_u2_u4_9254_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	142 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9254_Update/cr
      -- CP-element group 44: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9254_update_start_
      -- CP-element group 44: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9254_Update/$entry
      -- 
    cr_1259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(44), ack => CONCAT_u2_u4_9254_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	15 
    -- CP-element group 45: 	18 
    -- CP-element group 45: 	21 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9254_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9254_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9254_sample_completed_
      -- 
    ra_1255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u2_u4_9254_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	141 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9254_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9254_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9254_Update/ca
      -- 
    ca_1260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u2_u4_9254_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	142 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9258_update_start_
      -- CP-element group 47: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9258_Update/req
      -- CP-element group 47: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9258_Update/$entry
      -- 
    req_1273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(47), ack => W_issue_add_sub_9424_delayed_1_0_9256_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	20 
    -- CP-element group 48: successors 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	18 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9258_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9258_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9258_Sample/$exit
      -- 
    ack_1269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_issue_add_sub_9424_delayed_1_0_9256_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	141 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9258_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9258_Update/ack
      -- CP-element group 49: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9258_update_completed_
      -- 
    ack_1274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_issue_add_sub_9424_delayed_1_0_9256_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	17 
    -- CP-element group 50: 	20 
    -- CP-element group 50: 	23 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9266_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9266_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9266_Sample/$entry
      -- 
    rr_1282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(50), ack => CONCAT_u2_u4_9266_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	142 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9266_update_start_
      -- CP-element group 51: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9266_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9266_Update/cr
      -- 
    cr_1287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(51), ack => CONCAT_u2_u4_9266_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	15 
    -- CP-element group 52: 	18 
    -- CP-element group 52: 	21 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9266_Sample/ra
      -- CP-element group 52: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9266_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9266_sample_completed_
      -- 
    ra_1283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u2_u4_9266_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	141 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9266_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9266_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u2_u4_9266_Update/ca
      -- 
    ca_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u2_u4_9266_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	17 
    -- CP-element group 54: 	20 
    -- CP-element group 54: 	23 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9270_Sample/req
      -- CP-element group 54: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9270_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9270_sample_start_
      -- 
    req_1296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(54), ack => W_issue_div_9432_delayed_1_0_9268_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	142 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9270_update_start_
      -- CP-element group 55: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9270_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9270_Update/req
      -- 
    req_1301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(55), ack => W_issue_div_9432_delayed_1_0_9268_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	15 
    -- CP-element group 56: 	18 
    -- CP-element group 56: 	21 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9270_Sample/ack
      -- CP-element group 56: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9270_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9270_sample_completed_
      -- 
    ack_1297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_issue_div_9432_delayed_1_0_9268_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	141 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9270_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9270_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9270_Update/ack
      -- 
    ack_1302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_issue_div_9432_delayed_1_0_9268_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	17 
    -- CP-element group 58: 	20 
    -- CP-element group 58: 	23 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9296_start/req
      -- CP-element group 58: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9296_start/$entry
      -- CP-element group 58: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9296_sample_start_
      -- 
    req_1310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(58), ack => MUX_9296_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	142 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9296_complete/req
      -- CP-element group 59: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9296_complete/$entry
      -- CP-element group 59: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9296_update_start_
      -- 
    req_1315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(59), ack => MUX_9296_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	15 
    -- CP-element group 60: 	18 
    -- CP-element group 60: 	21 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9296_start/ack
      -- CP-element group 60: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9296_start/$exit
      -- CP-element group 60: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9296_sample_completed_
      -- 
    ack_1311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_9296_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	141 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9296_complete/ack
      -- CP-element group 61: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9296_complete/$exit
      -- CP-element group 61: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9296_update_completed_
      -- 
    ack_1316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_9296_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	17 
    -- CP-element group 62: 	23 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9318_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9318_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9318_Sample/rr
      -- 
    rr_1324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(62), ack => slice_9318_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	142 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9318_update_start_
      -- CP-element group 63: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9318_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9318_Update/cr
      -- 
    cr_1329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(63), ack => slice_9318_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	15 
    -- CP-element group 64: 	21 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9318_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9318_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9318_Sample/ra
      -- 
    ra_1325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_9318_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	141 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9318_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9318_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9318_Update/ca
      -- 
    ca_1330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_9318_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	17 
    -- CP-element group 66: 	23 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9322_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9322_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9322_Sample/rr
      -- 
    rr_1338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(66), ack => slice_9322_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	142 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9322_update_start_
      -- CP-element group 67: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9322_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9322_Update/cr
      -- 
    cr_1343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(67), ack => slice_9322_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	15 
    -- CP-element group 68: 	21 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9322_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9322_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9322_Sample/ra
      -- 
    ra_1339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_9322_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	141 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9322_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9322_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/slice_9322_Update/ca
      -- 
    ca_1344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_9322_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	142 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9333_update_start_
      -- CP-element group 70: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9333_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9333_Update/req
      -- 
    req_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(70), ack => W_issue_mul_9479_delayed_1_0_9331_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	20 
    -- CP-element group 71: successors 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	18 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9333_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9333_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9333_Sample/ack
      -- 
    ack_1353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_issue_mul_9479_delayed_1_0_9331_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	141 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9333_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9333_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9333_Update/ack
      -- 
    ack_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_issue_mul_9479_delayed_1_0_9331_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	17 
    -- CP-element group 73: 	20 
    -- CP-element group 73: 	23 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9336_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9336_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9336_Sample/req
      -- 
    req_1366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(73), ack => W_i32_mul_result_9480_delayed_1_0_9334_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	142 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9336_update_start_
      -- CP-element group 74: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9336_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9336_Update/req
      -- 
    req_1371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(74), ack => W_i32_mul_result_9480_delayed_1_0_9334_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	15 
    -- CP-element group 75: 	18 
    -- CP-element group 75: 	21 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9336_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9336_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9336_Sample/ack
      -- 
    ack_1367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_i32_mul_result_9480_delayed_1_0_9334_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	141 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9336_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9336_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9336_Update/ack
      -- 
    ack_1372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_i32_mul_result_9480_delayed_1_0_9334_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	17 
    -- CP-element group 77: 	20 
    -- CP-element group 77: 	23 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9347_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9347_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9347_start/req
      -- 
    req_1380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(77), ack => MUX_9347_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	142 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9347_update_start_
      -- CP-element group 78: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9347_complete/$entry
      -- CP-element group 78: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9347_complete/req
      -- 
    req_1385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(78), ack => MUX_9347_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	15 
    -- CP-element group 79: 	18 
    -- CP-element group 79: 	21 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9347_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9347_start/$exit
      -- CP-element group 79: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9347_start/ack
      -- 
    ack_1381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_9347_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	141 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9347_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9347_complete/$exit
      -- CP-element group 80: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/MUX_9347_complete/ack
      -- 
    ack_1386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_9347_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	17 
    -- CP-element group 81: 	20 
    -- CP-element group 81: 	23 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9351_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9351_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9351_Sample/req
      -- 
    req_1394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(81), ack => W_issue_div_9491_delayed_1_0_9349_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	142 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9351_update_start_
      -- CP-element group 82: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9351_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9351_Update/req
      -- 
    req_1399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(82), ack => W_issue_div_9491_delayed_1_0_9349_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	15 
    -- CP-element group 83: 	18 
    -- CP-element group 83: 	21 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9351_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9351_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9351_Sample/ack
      -- 
    ack_1395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_issue_div_9491_delayed_1_0_9349_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	141 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9351_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9351_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9351_Update/ack
      -- 
    ack_1400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_issue_div_9491_delayed_1_0_9349_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	17 
    -- CP-element group 85: 	20 
    -- CP-element group 85: 	23 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9361_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9361_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9361_Sample/rr
      -- 
    rr_1408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(85), ack => OR_u32_u32_9361_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	142 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9361_update_start_
      -- CP-element group 86: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9361_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9361_Update/cr
      -- 
    cr_1413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(86), ack => OR_u32_u32_9361_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	15 
    -- CP-element group 87: 	18 
    -- CP-element group 87: 	21 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9361_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9361_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9361_Sample/ra
      -- 
    ra_1409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_9361_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	141 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9361_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9361_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9361_Update/ca
      -- 
    ca_1414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_9361_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	17 
    -- CP-element group 89: 	20 
    -- CP-element group 89: 	23 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9382_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9382_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9382_Sample/rr
      -- 
    rr_1422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(89), ack => OR_u32_u32_9382_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	142 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9382_update_start_
      -- CP-element group 90: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9382_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9382_Update/cr
      -- 
    cr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(90), ack => OR_u32_u32_9382_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	15 
    -- CP-element group 91: 	18 
    -- CP-element group 91: 	21 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9382_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9382_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9382_Sample/ra
      -- 
    ra_1423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_9382_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	141 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9382_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9382_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u32_u32_9382_Update/ca
      -- 
    ca_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_9382_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	17 
    -- CP-element group 93: 	20 
    -- CP-element group 93: 	23 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9437_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9437_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9437_Sample/rr
      -- 
    rr_1436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(93), ack => OR_u1_u1_9437_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	142 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9437_update_start_
      -- CP-element group 94: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9437_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9437_Update/cr
      -- 
    cr_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(94), ack => OR_u1_u1_9437_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	15 
    -- CP-element group 95: 	18 
    -- CP-element group 95: 	21 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9437_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9437_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9437_Sample/ra
      -- 
    ra_1437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u1_u1_9437_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	141 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9437_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9437_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9437_Update/ca
      -- 
    ca_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u1_u1_9437_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	17 
    -- CP-element group 97: 	23 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9441_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9441_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9441_Sample/req
      -- 
    req_1450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(97), ack => W_psr_9567_delayed_1_0_9439_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	142 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9441_update_start_
      -- CP-element group 98: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9441_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9441_Update/req
      -- 
    req_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(98), ack => W_psr_9567_delayed_1_0_9439_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "iu_exec_daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	15 
    -- CP-element group 99: 	21 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9441_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9441_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9441_Sample/ack
      -- 
    ack_1451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_psr_9567_delayed_1_0_9439_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	141 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9441_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9441_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9441_Update/ack
      -- 
    ack_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_psr_9567_delayed_1_0_9439_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	142 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9444_update_start_
      -- CP-element group 101: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9444_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9444_Update/req
      -- 
    req_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(101), ack => W_exec_rett_9568_delayed_1_0_9442_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	20 
    -- CP-element group 102: successors 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	18 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9444_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9444_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9444_Sample/ack
      -- 
    ack_1465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_exec_rett_9568_delayed_1_0_9442_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	141 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9444_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9444_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9444_Update/ack
      -- 
    ack_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_exec_rett_9568_delayed_1_0_9442_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	17 
    -- CP-element group 104: 	20 
    -- CP-element group 104: 	23 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9447_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9447_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9447_Sample/req
      -- 
    req_1478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(104), ack => W_cti_next_psr_9569_delayed_1_0_9445_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	142 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9447_update_start_
      -- CP-element group 105: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9447_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9447_Update/req
      -- 
    req_1483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(105), ack => W_cti_next_psr_9569_delayed_1_0_9445_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	15 
    -- CP-element group 106: 	18 
    -- CP-element group 106: 	21 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9447_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9447_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9447_Sample/ack
      -- 
    ack_1479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_cti_next_psr_9569_delayed_1_0_9445_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	141 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9447_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9447_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9447_Update/ack
      -- 
    ack_1484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_cti_next_psr_9569_delayed_1_0_9445_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	142 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9450_update_start_
      -- CP-element group 108: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9450_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9450_Update/req
      -- 
    req_1497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(108), ack => W_write_psr_9570_delayed_1_0_9448_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	20 
    -- CP-element group 109: successors 
    -- CP-element group 109: marked-successors 
    -- CP-element group 109: 	18 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9450_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9450_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9450_Sample/ack
      -- 
    ack_1493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_psr_9570_delayed_1_0_9448_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	141 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9450_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9450_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9450_Update/ack
      -- 
    ack_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_psr_9570_delayed_1_0_9448_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	17 
    -- CP-element group 111: 	20 
    -- CP-element group 111: 	23 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9453_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9453_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9453_Sample/req
      -- 
    req_1506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(111), ack => W_i32_xor_result_9571_delayed_1_0_9451_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	142 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9453_update_start_
      -- CP-element group 112: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9453_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9453_Update/req
      -- 
    req_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(112), ack => W_i32_xor_result_9571_delayed_1_0_9451_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	15 
    -- CP-element group 113: 	18 
    -- CP-element group 113: 	21 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9453_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9453_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9453_Sample/ack
      -- 
    ack_1507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_i32_xor_result_9571_delayed_1_0_9451_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	141 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9453_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9453_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9453_Update/ack
      -- 
    ack_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_i32_xor_result_9571_delayed_1_0_9451_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	17 
    -- CP-element group 115: 	20 
    -- CP-element group 115: 	23 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9465_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9465_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9465_Sample/rr
      -- 
    rr_1520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(115), ack => OR_u1_u1_9465_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	142 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9465_update_start_
      -- CP-element group 116: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9465_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9465_Update/cr
      -- 
    cr_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(116), ack => OR_u1_u1_9465_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	15 
    -- CP-element group 117: 	18 
    -- CP-element group 117: 	21 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9465_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9465_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9465_Sample/ra
      -- 
    ra_1521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u1_u1_9465_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	141 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9465_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9465_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/OR_u1_u1_9465_Update/ca
      -- 
    ca_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u1_u1_9465_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	17 
    -- CP-element group 119: 	23 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9469_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9469_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9469_Sample/req
      -- 
    req_1534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(119), ack => W_psr_9584_delayed_1_0_9467_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	142 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9469_update_start_
      -- CP-element group 120: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9469_Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9469_Update/req
      -- 
    req_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(120), ack => W_psr_9584_delayed_1_0_9467_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	15 
    -- CP-element group 121: 	21 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9469_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9469_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9469_Sample/ack
      -- 
    ack_1535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_psr_9584_delayed_1_0_9467_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	141 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9469_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9469_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9469_Update/ack
      -- 
    ack_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_psr_9584_delayed_1_0_9467_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	17 
    -- CP-element group 123: 	20 
    -- CP-element group 123: 	23 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	125 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_to_stream_corrector_9734_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_to_stream_corrector_9734_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_to_stream_corrector_9734_Sample/req
      -- 
    req_1548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(123), ack => WPIPE_teu_iunit_to_stream_corrector_9734_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23) & iu_exec_daemon_CP_1081_elements(125);
      gj_iu_exec_daemon_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124: marked-successors 
    -- CP-element group 124: 	15 
    -- CP-element group 124: 	18 
    -- CP-element group 124: 	21 
    -- CP-element group 124:  members (6) 
      -- CP-element group 124: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_to_stream_corrector_9734_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_to_stream_corrector_9734_update_start_
      -- CP-element group 124: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_to_stream_corrector_9734_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_to_stream_corrector_9734_Sample/ack
      -- CP-element group 124: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_to_stream_corrector_9734_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_to_stream_corrector_9734_Update/req
      -- 
    ack_1549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_teu_iunit_to_stream_corrector_9734_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(124)); -- 
    req_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(124), ack => WPIPE_teu_iunit_to_stream_corrector_9734_inst_req_1); -- 
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	151 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	123 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_to_stream_corrector_9734_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_to_stream_corrector_9734_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_to_stream_corrector_9734_Update/ack
      -- 
    ack_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_teu_iunit_to_stream_corrector_9734_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	17 
    -- CP-element group 126: 	20 
    -- CP-element group 126: 	23 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u12_u14_9763_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u12_u14_9763_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u12_u14_9763_Sample/rr
      -- 
    rr_1562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(126), ack => CONCAT_u12_u14_9763_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	142 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u12_u14_9763_update_start_
      -- CP-element group 127: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u12_u14_9763_Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u12_u14_9763_Update/cr
      -- 
    cr_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(127), ack => CONCAT_u12_u14_9763_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: marked-successors 
    -- CP-element group 128: 	15 
    -- CP-element group 128: 	18 
    -- CP-element group 128: 	21 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u12_u14_9763_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u12_u14_9763_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u12_u14_9763_Sample/ra
      -- 
    ra_1563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u12_u14_9763_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	141 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u12_u14_9763_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u12_u14_9763_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u12_u14_9763_Update/ca
      -- 
    ca_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u12_u14_9763_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(129)); -- 
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	17 
    -- CP-element group 130: 	20 
    -- CP-element group 130: 	23 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u15_u16_9768_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u15_u16_9768_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u15_u16_9768_Sample/rr
      -- 
    rr_1576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(130), ack => CONCAT_u15_u16_9768_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	142 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u15_u16_9768_update_start_
      -- CP-element group 131: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u15_u16_9768_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u15_u16_9768_Update/cr
      -- 
    cr_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(131), ack => CONCAT_u15_u16_9768_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: marked-successors 
    -- CP-element group 132: 	15 
    -- CP-element group 132: 	18 
    -- CP-element group 132: 	21 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u15_u16_9768_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u15_u16_9768_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u15_u16_9768_Sample/ra
      -- 
    ra_1577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u15_u16_9768_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	141 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u15_u16_9768_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u15_u16_9768_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/CONCAT_u15_u16_9768_Update/ca
      -- 
    ca_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u15_u16_9768_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(133)); -- 
    -- CP-element group 134:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	17 
    -- CP-element group 134: 	20 
    -- CP-element group 134: 	23 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9772_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9772_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9772_Sample/req
      -- 
    req_1590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(134), ack => W_updated_y_9874_delayed_1_0_9770_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23);
      gj_iu_exec_daemon_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	142 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9772_update_start_
      -- CP-element group 135: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9772_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9772_Update/req
      -- 
    req_1595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(135), ack => W_updated_y_9874_delayed_1_0_9770_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: marked-successors 
    -- CP-element group 136: 	15 
    -- CP-element group 136: 	18 
    -- CP-element group 136: 	21 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9772_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9772_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9772_Sample/ack
      -- 
    ack_1591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_updated_y_9874_delayed_1_0_9770_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	141 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9772_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9772_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9772_Update/ack
      -- 
    ack_1596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_updated_y_9874_delayed_1_0_9770_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(137)); -- 
    -- CP-element group 138:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	142 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9786_update_start_
      -- CP-element group 138: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9786_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9786_Update/req
      -- 
    req_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(138), ack => W_send_to_wb_9880_delayed_1_0_9784_inst_req_1); -- 
    iu_exec_daemon_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= iu_exec_daemon_CP_1081_elements(142);
      gj_iu_exec_daemon_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	20 
    -- CP-element group 139: successors 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	18 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9786_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9786_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9786_Sample/ack
      -- 
    ack_1605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_to_wb_9880_delayed_1_0_9784_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9786_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9786_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/assign_stmt_9786_Update/ack
      -- 
    ack_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_to_wb_9880_delayed_1_0_9784_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(140)); -- 
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	96 
    -- CP-element group 141: 	76 
    -- CP-element group 141: 	80 
    -- CP-element group 141: 	84 
    -- CP-element group 141: 	69 
    -- CP-element group 141: 	88 
    -- CP-element group 141: 	92 
    -- CP-element group 141: 	118 
    -- CP-element group 141: 	122 
    -- CP-element group 141: 	129 
    -- CP-element group 141: 	133 
    -- CP-element group 141: 	137 
    -- CP-element group 141: 	140 
    -- CP-element group 141: 	72 
    -- CP-element group 141: 	110 
    -- CP-element group 141: 	114 
    -- CP-element group 141: 	103 
    -- CP-element group 141: 	107 
    -- CP-element group 141: 	100 
    -- CP-element group 141: 	39 
    -- CP-element group 141: 	42 
    -- CP-element group 141: 	46 
    -- CP-element group 141: 	49 
    -- CP-element group 141: 	53 
    -- CP-element group 141: 	57 
    -- CP-element group 141: 	61 
    -- CP-element group 141: 	65 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_to_writeback_9788_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_to_writeback_9788_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_to_writeback_9788_Sample/req
      -- 
    req_1618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(141), ack => WPIPE_iunit_exec_to_writeback_9788_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 27) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1);
      constant place_markings: IntegerArray(0 to 27)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 1);
      constant place_delays: IntegerArray(0 to 27) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 28); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(96) & iu_exec_daemon_CP_1081_elements(76) & iu_exec_daemon_CP_1081_elements(80) & iu_exec_daemon_CP_1081_elements(84) & iu_exec_daemon_CP_1081_elements(69) & iu_exec_daemon_CP_1081_elements(88) & iu_exec_daemon_CP_1081_elements(92) & iu_exec_daemon_CP_1081_elements(118) & iu_exec_daemon_CP_1081_elements(122) & iu_exec_daemon_CP_1081_elements(129) & iu_exec_daemon_CP_1081_elements(133) & iu_exec_daemon_CP_1081_elements(137) & iu_exec_daemon_CP_1081_elements(140) & iu_exec_daemon_CP_1081_elements(72) & iu_exec_daemon_CP_1081_elements(110) & iu_exec_daemon_CP_1081_elements(114) & iu_exec_daemon_CP_1081_elements(103) & iu_exec_daemon_CP_1081_elements(107) & iu_exec_daemon_CP_1081_elements(100) & iu_exec_daemon_CP_1081_elements(39) & iu_exec_daemon_CP_1081_elements(42) & iu_exec_daemon_CP_1081_elements(46) & iu_exec_daemon_CP_1081_elements(49) & iu_exec_daemon_CP_1081_elements(53) & iu_exec_daemon_CP_1081_elements(57) & iu_exec_daemon_CP_1081_elements(61) & iu_exec_daemon_CP_1081_elements(65) & iu_exec_daemon_CP_1081_elements(143);
      gj_iu_exec_daemon_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 28, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	94 
    -- CP-element group 142: 	74 
    -- CP-element group 142: 	90 
    -- CP-element group 142: 	82 
    -- CP-element group 142: 	86 
    -- CP-element group 142: 	78 
    -- CP-element group 142: 	70 
    -- CP-element group 142: 	120 
    -- CP-element group 142: 	127 
    -- CP-element group 142: 	131 
    -- CP-element group 142: 	135 
    -- CP-element group 142: 	138 
    -- CP-element group 142: 	112 
    -- CP-element group 142: 	116 
    -- CP-element group 142: 	105 
    -- CP-element group 142: 	108 
    -- CP-element group 142: 	98 
    -- CP-element group 142: 	101 
    -- CP-element group 142: 	37 
    -- CP-element group 142: 	40 
    -- CP-element group 142: 	44 
    -- CP-element group 142: 	47 
    -- CP-element group 142: 	51 
    -- CP-element group 142: 	55 
    -- CP-element group 142: 	59 
    -- CP-element group 142: 	63 
    -- CP-element group 142: 	67 
    -- CP-element group 142:  members (6) 
      -- CP-element group 142: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_to_writeback_9788_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_to_writeback_9788_update_start_
      -- CP-element group 142: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_to_writeback_9788_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_to_writeback_9788_Sample/ack
      -- CP-element group 142: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_to_writeback_9788_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_to_writeback_9788_Update/req
      -- 
    ack_1619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_iunit_exec_to_writeback_9788_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(142)); -- 
    req_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(142), ack => WPIPE_iunit_exec_to_writeback_9788_inst_req_1); -- 
    -- CP-element group 143:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	151 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_to_writeback_9788_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_to_writeback_9788_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_iunit_exec_to_writeback_9788_Update/ack
      -- 
    ack_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_iunit_exec_to_writeback_9788_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(143)); -- 
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	17 
    -- CP-element group 144: 	20 
    -- CP-element group 144: 	23 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_loadstore_9821_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_loadstore_9821_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_loadstore_9821_Sample/req
      -- 
    req_1632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(144), ack => WPIPE_teu_iunit_trap_to_loadstore_9821_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23) & iu_exec_daemon_CP_1081_elements(146);
      gj_iu_exec_daemon_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	15 
    -- CP-element group 145: 	18 
    -- CP-element group 145: 	21 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_loadstore_9821_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_loadstore_9821_update_start_
      -- CP-element group 145: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_loadstore_9821_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_loadstore_9821_Sample/ack
      -- CP-element group 145: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_loadstore_9821_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_loadstore_9821_Update/req
      -- 
    ack_1633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_teu_iunit_trap_to_loadstore_9821_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(145)); -- 
    req_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(145), ack => WPIPE_teu_iunit_trap_to_loadstore_9821_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	151 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_loadstore_9821_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_loadstore_9821_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_loadstore_9821_Update/ack
      -- 
    ack_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_teu_iunit_trap_to_loadstore_9821_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	17 
    -- CP-element group 147: 	20 
    -- CP-element group 147: 	23 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_fpunit_9840_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_fpunit_9840_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_fpunit_9840_Sample/req
      -- 
    req_1646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(147), ack => WPIPE_teu_iunit_trap_to_fpunit_9840_inst_req_0); -- 
    iu_exec_daemon_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(17) & iu_exec_daemon_CP_1081_elements(20) & iu_exec_daemon_CP_1081_elements(23) & iu_exec_daemon_CP_1081_elements(149);
      gj_iu_exec_daemon_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	15 
    -- CP-element group 148: 	18 
    -- CP-element group 148: 	21 
    -- CP-element group 148:  members (6) 
      -- CP-element group 148: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_fpunit_9840_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_fpunit_9840_update_start_
      -- CP-element group 148: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_fpunit_9840_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_fpunit_9840_Sample/ack
      -- CP-element group 148: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_fpunit_9840_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_fpunit_9840_Update/req
      -- 
    ack_1647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_teu_iunit_trap_to_fpunit_9840_inst_ack_0, ack => iu_exec_daemon_CP_1081_elements(148)); -- 
    req_1651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(148), ack => WPIPE_teu_iunit_trap_to_fpunit_9840_inst_req_1); -- 
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	147 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_fpunit_9840_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_fpunit_9840_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/WPIPE_teu_iunit_trap_to_fpunit_9840_Update/ack
      -- 
    ack_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_teu_iunit_trap_to_fpunit_9840_inst_ack_1, ack => iu_exec_daemon_CP_1081_elements(149)); -- 
    -- CP-element group 150:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	9 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	5 
    -- CP-element group 150:  members (2) 
      -- CP-element group 150: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/condition_evaluated
      -- CP-element group 150: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/loop_body_delay_to_condition_start
      -- 
    condition_evaluated_1105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => iu_exec_daemon_CP_1081_elements(150), ack => do_while_stmt_8361_branch_req_0); -- 
    -- Element group iu_exec_daemon_CP_1081_elements(150) is a control-delay.
    cp_element_150_delay: control_delay_element  generic map(name => " 150_delay", delay_value => 1)  port map(req => iu_exec_daemon_CP_1081_elements(9), ack => iu_exec_daemon_CP_1081_elements(150), clk => clk, reset =>reset);
    -- CP-element group 151:  join  transition  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	125 
    -- CP-element group 151: 	143 
    -- CP-element group 151: 	146 
    -- CP-element group 151: 	149 
    -- CP-element group 151: 	26 
    -- CP-element group 151: 	29 
    -- CP-element group 151: 	32 
    -- CP-element group 151: 	35 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	6 
    -- CP-element group 151:  members (1) 
      -- CP-element group 151: 	 branch_block_stmt_8360/do_while_stmt_8361/do_while_stmt_8361_loop_body/$exit
      -- 
    iu_exec_daemon_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 7);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 35) := "iu_exec_daemon_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= iu_exec_daemon_CP_1081_elements(125) & iu_exec_daemon_CP_1081_elements(143) & iu_exec_daemon_CP_1081_elements(146) & iu_exec_daemon_CP_1081_elements(149) & iu_exec_daemon_CP_1081_elements(26) & iu_exec_daemon_CP_1081_elements(29) & iu_exec_daemon_CP_1081_elements(32) & iu_exec_daemon_CP_1081_elements(35);
      gj_iu_exec_daemon_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	5 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (2) 
      -- CP-element group 152: 	 branch_block_stmt_8360/do_while_stmt_8361/loop_exit/$exit
      -- CP-element group 152: 	 branch_block_stmt_8360/do_while_stmt_8361/loop_exit/ack
      -- 
    ack_1657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_8361_branch_ack_0, ack => iu_exec_daemon_CP_1081_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	5 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (2) 
      -- CP-element group 153: 	 branch_block_stmt_8360/do_while_stmt_8361/loop_taken/$exit
      -- CP-element group 153: 	 branch_block_stmt_8360/do_while_stmt_8361/loop_taken/ack
      -- 
    ack_1661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_8361_branch_ack_1, ack => iu_exec_daemon_CP_1081_elements(153)); -- 
    -- CP-element group 154:  transition  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	3 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	1 
    -- CP-element group 154:  members (1) 
      -- CP-element group 154: 	 branch_block_stmt_8360/do_while_stmt_8361/$exit
      -- 
    iu_exec_daemon_CP_1081_elements(154) <= iu_exec_daemon_CP_1081_elements(3);
    iu_exec_daemon_do_while_stmt_8361_terminator_1662: loop_terminator -- 
      generic map (name => " iu_exec_daemon_do_while_stmt_8361_terminator_1662", max_iterations_in_flight =>7) 
      port map(loop_body_exit => iu_exec_daemon_CP_1081_elements(6),loop_continue => iu_exec_daemon_CP_1081_elements(153),loop_terminate => iu_exec_daemon_CP_1081_elements(152),loop_back => iu_exec_daemon_CP_1081_elements(4),loop_exit => iu_exec_daemon_CP_1081_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_1106_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= iu_exec_daemon_CP_1081_elements(7);
        preds(1)  <= iu_exec_daemon_CP_1081_elements(8);
        entry_tmerge_1106 : transition_merge -- 
          generic map(name => " entry_tmerge_1106")
          port map (preds => preds, symbol_out => iu_exec_daemon_CP_1081_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_9066_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9073_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9083_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9090_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9110_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9197_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9207_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9240_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9464_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9493_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9501_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9540_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9553_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9566_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9589_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9592_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9616_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9680_wire : std_logic_vector(0 downto 0);
    signal AND_u32_u32_8756_wire : std_logic_vector(31 downto 0);
    signal BITSEL_u32_u1_8783_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_9492_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_9504_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u12_u14_9868_9868_delayed_1_0_9764 : std_logic_vector(13 downto 0);
    signal CONCAT_u12_u32_9102_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u13_u20_9715_wire : std_logic_vector(19 downto 0);
    signal CONCAT_u15_u16_9871_9871_delayed_1_0_9769 : std_logic_vector(15 downto 0);
    signal CONCAT_u16_u48_9777_wire : std_logic_vector(47 downto 0);
    signal CONCAT_u1_u2_9029_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9032_wire_constant : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9037_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9040_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9045_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9048_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9052_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9055_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9250_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9253_wire_constant : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9262_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9265_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9275_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9278_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9283_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9286_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9290_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9293_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9306_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9309_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9642_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9647_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9651_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9710_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9718_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9721_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9725_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9762_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u5_9117_wire : std_logic_vector(4 downto 0);
    signal CONCAT_u1_u5_9149_wire : std_logic_vector(4 downto 0);
    signal CONCAT_u1_u5_9713_wire : std_logic_vector(4 downto 0);
    signal CONCAT_u1_u6_9124_wire : std_logic_vector(5 downto 0);
    signal CONCAT_u1_u8_9654_wire : std_logic_vector(7 downto 0);
    signal CONCAT_u2_u10_9655_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u2_u3_9644_wire : std_logic_vector(2 downto 0);
    signal CONCAT_u2_u4_9033_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_9041_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_9049_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_9056_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_9279_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_9287_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_9294_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_9310_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_9423_9423_delayed_1_0_9255 : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_9431_9431_delayed_1_0_9267 : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_9722_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u66_9729_wire : std_logic_vector(65 downto 0);
    signal CONCAT_u2_u7_9714_wire : std_logic_vector(6 downto 0);
    signal CONCAT_u2_u8_9120_wire : std_logic_vector(7 downto 0);
    signal CONCAT_u32_u64_9127_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_9176_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_9728_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_9780_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u3_u5_9648_wire : std_logic_vector(4 downto 0);
    signal CONCAT_u48_u112_9781_wire : std_logic_vector(111 downto 0);
    signal CONCAT_u4_u6_9169_wire : std_logic_vector(5 downto 0);
    signal CONCAT_u4_u6_9703_wire : std_logic_vector(5 downto 0);
    signal CONCAT_u4_u6_9757_wire : std_logic_vector(5 downto 0);
    signal CONCAT_u4_u6_9833_wire : std_logic_vector(5 downto 0);
    signal CONCAT_u4_u70_9730_wire : std_logic_vector(69 downto 0);
    signal CONCAT_u5_u13_9121_wire : std_logic_vector(12 downto 0);
    signal CONCAT_u5_u7_9151_wire : std_logic_vector(6 downto 0);
    signal CONCAT_u64_u96_9178_wire : std_logic_vector(95 downto 0);
    signal CONCAT_u6_u10_9154_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u6_u12_9759_wire : std_logic_vector(11 downto 0);
    signal CONCAT_u6_u13_9173_wire : std_logic_vector(12 downto 0);
    signal CONCAT_u6_u13_9707_wire : std_logic_vector(12 downto 0);
    signal CONCAT_u6_u70_9128_wire : std_logic_vector(69 downto 0);
    signal CONCAT_u6_u7_9172_wire : std_logic_vector(6 downto 0);
    signal CONCAT_u6_u7_9706_wire : std_logic_vector(6 downto 0);
    signal CONCAT_u6_u7_9836_wire : std_logic_vector(6 downto 0);
    signal CONCAT_u8_u12_9099_wire : std_logic_vector(11 downto 0);
    signal CONCAT_u8_u12_9327_wire : std_logic_vector(11 downto 0);
    signal Caddsub_8727 : std_logic_vector(0 downto 0);
    signal Cdiv_9223 : std_logic_vector(0 downto 0);
    signal Ci_8697 : std_logic_vector(0 downto 0);
    signal Clogical_8806 : std_logic_vector(0 downto 0);
    signal Cmul_8878 : std_logic_vector(0 downto 0);
    signal Cmulscc_8843 : std_logic_vector(0 downto 0);
    signal EQ_u32_u1_8791_wire : std_logic_vector(0 downto 0);
    signal EQ_u32_u1_9200_wire : std_logic_vector(0 downto 0);
    signal MUX_8758_wire : std_logic_vector(31 downto 0);
    signal MUX_8764_wire : std_logic_vector(31 downto 0);
    signal MUX_8769_wire : std_logic_vector(31 downto 0);
    signal MUX_8775_wire : std_logic_vector(31 downto 0);
    signal MUX_8995_wire : std_logic_vector(31 downto 0);
    signal MUX_9002_wire : std_logic_vector(31 downto 0);
    signal MUX_9006_wire : std_logic_vector(31 downto 0);
    signal MUX_9011_wire : std_logic_vector(31 downto 0);
    signal MUX_9015_wire : std_logic_vector(31 downto 0);
    signal MUX_9057_wire : std_logic_vector(3 downto 0);
    signal MUX_9058_wire : std_logic_vector(3 downto 0);
    signal MUX_9295_wire : std_logic_vector(3 downto 0);
    signal MUX_9312_wire : std_logic_vector(3 downto 0);
    signal MUX_9313_wire : std_logic_vector(3 downto 0);
    signal MUX_9356_wire : std_logic_vector(31 downto 0);
    signal MUX_9360_wire : std_logic_vector(31 downto 0);
    signal MUX_9367_wire : std_logic_vector(31 downto 0);
    signal MUX_9371_wire : std_logic_vector(31 downto 0);
    signal MUX_9376_wire : std_logic_vector(31 downto 0);
    signal MUX_9380_wire : std_logic_vector(31 downto 0);
    signal MUX_9391_wire : std_logic_vector(31 downto 0);
    signal MUX_9464_9464_delayed_1_0_9297 : std_logic_vector(3 downto 0);
    signal MUX_9480_wire : std_logic_vector(31 downto 0);
    signal MUX_9481_wire : std_logic_vector(31 downto 0);
    signal MUX_9482_wire : std_logic_vector(31 downto 0);
    signal MUX_9490_9490_delayed_1_0_9348 : std_logic_vector(31 downto 0);
    signal MUX_9549_wire : std_logic_vector(31 downto 0);
    signal MUX_9556_wire : std_logic_vector(31 downto 0);
    signal MUX_9625_wire : std_logic_vector(0 downto 0);
    signal MUX_9629_wire : std_logic_vector(0 downto 0);
    signal NEQ_u6_u1_9683_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8609_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8614_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8620_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8626_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8632_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8638_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8644_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8700_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8730_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8809_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8826_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8846_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8896_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8902_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8908_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8914_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8920_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8926_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_8983_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9063_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9065_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9080_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9082_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9107_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9109_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9195_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9205_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9209_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9487_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9499_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9505_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9510_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9520_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9533_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9551_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9562_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9585_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9588_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9613_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9621_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_9677_wire : std_logic_vector(0 downto 0);
    signal NOT_u32_u32_8743_wire : std_logic_vector(31 downto 0);
    signal Naddsub_8727 : std_logic_vector(0 downto 0);
    signal Ndiv_9223 : std_logic_vector(0 downto 0);
    signal Ni_8682 : std_logic_vector(0 downto 0);
    signal Nlogical_8786 : std_logic_vector(0 downto 0);
    signal Nmul_8867 : std_logic_vector(0 downto 0);
    signal Nmulscc_8843 : std_logic_vector(0 downto 0);
    signal OR_u1_u1_8663_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_8666_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_8667_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_8703_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_8733_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_8736_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_8737_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_8812_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_8814_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_8986_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9069_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9071_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9075_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9087_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9089_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9227_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9229_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9232_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9234_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9340_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9343_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9344_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9459_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9462_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9463_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9494_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9523_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9566_9566_delayed_1_0_9438 : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9567_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9582_9582_delayed_1_0_9466 : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9593_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9630_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9661_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9664_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9665_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9668_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9671_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9672_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9684_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_8762_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_8765_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_8776_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_9007_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_9016_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_9372_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_9381_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_9392_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_9394_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_9396_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_9504_9504_delayed_1_0_9362 : std_logic_vector(31 downto 0);
    signal OR_u32_u32_9524_9524_delayed_1_0_9383 : std_logic_vector(31 downto 0);
    signal OR_u32_u32_9557_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_8534_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_7_9636_wire_constant : std_logic_vector(6 downto 0);
    signal S_9582 : std_logic_vector(0 downto 0);
    signal UGE_u5_u1_9539_wire : std_logic_vector(0 downto 0);
    signal Vaddsub_8727 : std_logic_vector(0 downto 0);
    signal Vdiv_9223 : std_logic_vector(0 downto 0);
    signal Vi_8692 : std_logic_vector(0 downto 0);
    signal Vlogical_8800 : std_logic_vector(0 downto 0);
    signal Vmul_8875 : std_logic_vector(0 downto 0);
    signal Vmulscc_8843 : std_logic_vector(0 downto 0);
    signal XOR_u32_u32_8773_wire : std_logic_vector(31 downto 0);
    signal Zaddsub_8727 : std_logic_vector(0 downto 0);
    signal Zdiv_9223 : std_logic_vector(0 downto 0);
    signal Zi_8687 : std_logic_vector(0 downto 0);
    signal Zlogical_8794 : std_logic_vector(0 downto 0);
    signal Zmul_8872 : std_logic_vector(0 downto 0);
    signal Zmulscc_8843 : std_logic_vector(0 downto 0);
    signal alu_8605 : std_logic_vector(0 downto 0);
    signal alu_cc_flags_9315 : std_logic_vector(3 downto 0);
    signal alu_overflow_trap_9600 : std_logic_vector(0 downto 0);
    signal alu_psr_9330 : std_logic_vector(31 downto 0);
    signal alu_result_9398 : std_logic_vector(31 downto 0);
    signal alu_trap_9243 : std_logic_vector(0 downto 0);
    signal alu_was_used_9236 : std_logic_vector(0 downto 0);
    signal annul_flag_8605 : std_logic_vector(0 downto 0);
    signal annul_next_9696 : std_logic_vector(0 downto 0);
    signal asr_8547 : std_logic_vector(31 downto 0);
    signal asr_id_8605 : std_logic_vector(4 downto 0);
    signal br_cond_8605 : std_logic_vector(3 downto 0);
    signal br_taken_9691 : std_logic_vector(0 downto 0);
    signal bypass_cc_to_reg_file_9156 : std_logic_vector(16 downto 0);
    signal bypass_to_reg_file_9130 : std_logic_vector(82 downto 0);
    signal cti_8605 : std_logic_vector(0 downto 0);
    signal cti_annul_next_8951 : std_logic_vector(0 downto 0);
    signal cti_br_taken_8951 : std_logic_vector(0 downto 0);
    signal cti_illegal_instr_trap_8951 : std_logic_vector(0 downto 0);
    signal cti_mem_address_not_aligned_trap_8951 : std_logic_vector(0 downto 0);
    signal cti_next_psr_8951 : std_logic_vector(31 downto 0);
    signal cti_next_psr_9569_delayed_1_0_9447 : std_logic_vector(31 downto 0);
    signal cti_privileged_instr_trap_8951 : std_logic_vector(0 downto 0);
    signal cti_processor_error_mode_8951 : std_logic_vector(0 downto 0);
    signal cti_ticc_trap_type_8951 : std_logic_vector(6 downto 0);
    signal cti_trap_8956 : std_logic_vector(0 downto 0);
    signal cti_trap_instr_trap_8951 : std_logic_vector(0 downto 0);
    signal cti_trap_status_8951 : std_logic_vector(0 downto 0);
    signal cti_window_underflow_trap_8951 : std_logic_vector(0 downto 0);
    signal div_by_0_trap_9202 : std_logic_vector(0 downto 0);
    signal do_not_bypass_8399 : std_logic_vector(0 downto 0);
    signal dti_8605 : std_logic_vector(0 downto 0);
    signal exec_bicc_8923 : std_logic_vector(0 downto 0);
    signal exec_call_8899 : std_logic_vector(0 downto 0);
    signal exec_control_word_8395 : std_logic_vector(54 downto 0);
    signal exec_info_8365 : std_logic_vector(149 downto 0);
    signal exec_info_d_8379 : std_logic_vector(149 downto 0);
    signal exec_jmpl_8911 : std_logic_vector(0 downto 0);
    signal exec_processor_error_mode_9686 : std_logic_vector(0 downto 0);
    signal exec_rett_8905 : std_logic_vector(0 downto 0);
    signal exec_rett_9568_delayed_1_0_9444 : std_logic_vector(0 downto 0);
    signal exec_ticc_8917 : std_logic_vector(0 downto 0);
    signal fast_alu_cc_flags_9060 : std_logic_vector(3 downto 0);
    signal fast_alu_psr_9104 : std_logic_vector(31 downto 0);
    signal fast_alu_result_9024 : std_logic_vector(31 downto 0);
    signal fast_fast_alu_result_9018 : std_logic_vector(31 downto 0);
    signal fast_result_to_wb_9180 : std_logic_vector(108 downto 0);
    signal fast_update_psr_9077 : std_logic_vector(0 downto 0);
    signal get_from_rfile_8370 : std_logic_vector(0 downto 0);
    signal get_from_rfile_8647_delayed_1_0_8478 : std_logic_vector(0 downto 0);
    signal i32_add_sub_ovflow_trap_8727 : std_logic_vector(0 downto 0);
    signal i32_add_sub_result_8727 : std_logic_vector(31 downto 0);
    signal i32_div_result_9223 : std_logic_vector(31 downto 0);
    signal i32_logical_op_result_8778 : std_logic_vector(31 downto 0);
    signal i32_mul_result_8857 : std_logic_vector(31 downto 0);
    signal i32_mul_result_9480_delayed_1_0_9336 : std_logic_vector(31 downto 0);
    signal i32_mul_y_8893 : std_logic_vector(31 downto 0);
    signal i32_mulscc_result_8843 : std_logic_vector(31 downto 0);
    signal i32_mulscc_y_8843 : std_logic_vector(31 downto 0);
    signal i32_shift_result_8823 : std_logic_vector(31 downto 0);
    signal i32_xor_result_8751 : std_logic_vector(31 downto 0);
    signal i32_xor_result_9571_delayed_1_0_9453 : std_logic_vector(31 downto 0);
    signal illegal_instr_trap_9569 : std_logic_vector(0 downto 0);
    signal imm_flag_8403 : std_logic_vector(0 downto 0);
    signal imm_operand_8451 : std_logic_vector(31 downto 0);
    signal is_bicc_8605 : std_logic_vector(0 downto 0);
    signal is_call_8605 : std_logic_vector(0 downto 0);
    signal is_cbccc_8605 : std_logic_vector(0 downto 0);
    signal is_fbfcc_8605 : std_logic_vector(0 downto 0);
    signal is_jmpl_8605 : std_logic_vector(0 downto 0);
    signal is_load_to_debug_8605 : std_logic_vector(0 downto 0);
    signal is_restore_8605 : std_logic_vector(0 downto 0);
    signal is_rett_8605 : std_logic_vector(0 downto 0);
    signal is_save_8605 : std_logic_vector(0 downto 0);
    signal is_sethi_8605 : std_logic_vector(0 downto 0);
    signal is_store_to_debug_8605 : std_logic_vector(0 downto 0);
    signal is_ticc_8605 : std_logic_vector(0 downto 0);
    signal issue_add_sub_8705 : std_logic_vector(0 downto 0);
    signal issue_add_sub_9424_delayed_1_0_9258 : std_logic_vector(0 downto 0);
    signal issue_cti_8929 : std_logic_vector(0 downto 0);
    signal issue_div_9211 : std_logic_vector(0 downto 0);
    signal issue_div_9432_delayed_1_0_9270 : std_logic_vector(0 downto 0);
    signal issue_div_9491_delayed_1_0_9351 : std_logic_vector(0 downto 0);
    signal issue_logical_8739 : std_logic_vector(0 downto 0);
    signal issue_mul_8849 : std_logic_vector(0 downto 0);
    signal issue_mul_9416_delayed_1_0_9246 : std_logic_vector(0 downto 0);
    signal issue_mul_9479_delayed_1_0_9333 : std_logic_vector(0 downto 0);
    signal issue_mulscc_8829 : std_logic_vector(0 downto 0);
    signal issue_read_asr_8647 : std_logic_vector(0 downto 0);
    signal issue_read_psr_8623 : std_logic_vector(0 downto 0);
    signal issue_read_tbr_8635 : std_logic_vector(0 downto 0);
    signal issue_read_wim_8629 : std_logic_vector(0 downto 0);
    signal issue_read_y_8641 : std_logic_vector(0 downto 0);
    signal issue_sethi_8617 : std_logic_vector(0 downto 0);
    signal issue_shift_8816 : std_logic_vector(0 downto 0);
    signal iu1_to_cu2_8443 : std_logic_vector(0 downto 0);
    signal iu1_to_fu2_8439 : std_logic_vector(0 downto 0);
    signal iu1_to_iu2_8423 : std_logic_vector(0 downto 0);
    signal iu1_to_ls_trap_8435 : std_logic_vector(0 downto 0);
    signal iu1_to_sc_8427 : std_logic_vector(0 downto 0);
    signal iu_S_9530 : std_logic_vector(0 downto 0);
    signal iu_disable_traps_9507 : std_logic_vector(0 downto 0);
    signal iu_dti_8605 : std_logic_vector(0 downto 0);
    signal iu_enable_traps_9496 : std_logic_vector(0 downto 0);
    signal iu_proc_ilvl_9517 : std_logic_vector(3 downto 0);
    signal iu_reg_to_ls_8431 : std_logic_vector(0 downto 0);
    signal iu_set_S_9525 : std_logic_vector(0 downto 0);
    signal iu_set_proc_ilvl_9513 : std_logic_vector(0 downto 0);
    signal iu_to_fu_trapped_9829 : std_logic_vector(0 downto 0);
    signal iu_to_ls_trapped_9819 : std_logic_vector(0 downto 0);
    signal iunit_has_trapped_9674 : std_logic_vector(0 downto 0);
    signal konst_8368_wire_constant : std_logic_vector(149 downto 0);
    signal konst_8482_wire_constant : std_logic_vector(141 downto 0);
    signal konst_8680_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8685_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8690_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8695_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8757_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8763_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8768_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8774_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8782_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8790_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8797_wire_constant : std_logic_vector(0 downto 0);
    signal konst_8803_wire_constant : std_logic_vector(0 downto 0);
    signal konst_8865_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8870_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8882_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9001_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9005_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9010_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9014_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9199_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9346_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9355_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9359_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9366_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9370_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9375_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9379_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9390_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9491_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9503_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9528_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9548_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9555_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9580_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9624_wire_constant : std_logic_vector(0 downto 0);
    signal konst_9628_wire_constant : std_logic_vector(0 downto 0);
    signal konst_9848_wire_constant : std_logic_vector(0 downto 0);
    signal l_operand_2_8746 : std_logic_vector(31 downto 0);
    signal mem_addr_not_aligned_trap_9610 : std_logic_vector(0 downto 0);
    signal misc_8605 : std_logic_vector(0 downto 0);
    signal mul_y_op_1_8884 : std_logic_vector(31 downto 0);
    signal mul_y_op_2_8888 : std_logic_vector(31 downto 0);
    signal negate_second_operand_8605 : std_logic_vector(0 downto 0);
    signal operand_1_8671 : std_logic_vector(31 downto 0);
    signal operand_2_8677 : std_logic_vector(31 downto 0);
    signal ops_8376 : std_logic_vector(141 downto 0);
    signal ops_qualified_8484 : std_logic_vector(141 downto 0);
    signal ops_valid_8492 : std_logic_vector(0 downto 0);
    signal pc_8455 : std_logic_vector(31 downto 0);
    signal post_rett_or_write_psr_psr_8997 : std_logic_vector(31 downto 0);
    signal priv_instr_trap_9595 : std_logic_vector(0 downto 0);
    signal psr_8516 : std_logic_vector(31 downto 0);
    signal psr_9567_delayed_1_0_9441 : std_logic_vector(31 downto 0);
    signal psr_9584_delayed_1_0_9469 : std_logic_vector(31 downto 0);
    signal rd_8411 : std_logic_vector(4 downto 0);
    signal read_asr_8605 : std_logic_vector(0 downto 0);
    signal read_psr_8605 : std_logic_vector(0 downto 0);
    signal read_tbr_8605 : std_logic_vector(0 downto 0);
    signal read_wim_8605 : std_logic_vector(0 downto 0);
    signal read_y_8605 : std_logic_vector(0 downto 0);
    signal restore_uflow_trap_8555 : std_logic_vector(0 downto 0);
    signal rf_operand_1_8508 : std_logic_vector(31 downto 0);
    signal rf_operand_2_8512 : std_logic_vector(31 downto 0);
    signal save_ovflow_trap_8551 : std_logic_vector(0 downto 0);
    signal send_alu_bypass_9113 : std_logic_vector(0 downto 0);
    signal send_cc_bypass_9092 : std_logic_vector(0 downto 0);
    signal send_fast_alu_result_8419 : std_logic_vector(0 downto 0);
    signal send_to_sc_9699 : std_logic_vector(0 downto 0);
    signal send_to_wb_9753 : std_logic_vector(0 downto 0);
    signal send_to_wb_9880_delayed_1_0_9786 : std_logic_vector(0 downto 0);
    signal set_cc_8605 : std_logic_vector(0 downto 0);
    signal signed_correction_8862 : std_logic_vector(31 downto 0);
    signal signed_mul_div_8605 : std_logic_vector(0 downto 0);
    signal skip_alu_exec_8611 : std_logic_vector(0 downto 0);
    signal skip_from_rfile_8488 : std_logic_vector(0 downto 0);
    signal skip_iu_8447 : std_logic_vector(0 downto 0);
    signal slice_9097_wire : std_logic_vector(7 downto 0);
    signal slice_9101_wire : std_logic_vector(19 downto 0);
    signal slice_9471_9471_delayed_1_0_9319 : std_logic_vector(7 downto 0);
    signal slice_9475_9475_delayed_1_0_9323 : std_logic_vector(19 downto 0);
    signal slice_9536_wire : std_logic_vector(4 downto 0);
    signal slot_id_1_8504 : std_logic_vector(5 downto 0);
    signal slot_id_8391 : std_logic_vector(5 downto 0);
    signal sr_illegal_instr_trap_9542 : std_logic_vector(0 downto 0);
    signal sreg_value_8520 : std_logic_vector(31 downto 0);
    signal stream_id_1_8500 : std_logic_vector(1 downto 0);
    signal stream_id_8387 : std_logic_vector(1 downto 0);
    signal tagged_alu_op_8605 : std_logic_vector(0 downto 0);
    signal tbr_8541 : std_logic_vector(31 downto 0);
    signal thread_id_1_8496 : std_logic_vector(3 downto 0);
    signal thread_id_8383 : std_logic_vector(3 downto 0);
    signal ticc_trap_type_9638 : std_logic_vector(6 downto 0);
    signal to_fpu_9838 : std_logic_vector(12 downto 0);
    signal to_iu_wb_9783 : std_logic_vector(125 downto 0);
    signal to_sc_9732 : std_logic_vector(89 downto 0);
    signal trap_if_not_super_8407 : std_logic_vector(0 downto 0);
    signal trap_instr_trap_9605 : std_logic_vector(0 downto 0);
    signal trap_on_overflow_8605 : std_logic_vector(0 downto 0);
    signal trap_or_error_9816 : std_logic_vector(0 downto 0);
    signal traps_9657 : std_logic_vector(14 downto 0);
    signal type_cast_9538_wire_constant : std_logic_vector(4 downto 0);
    signal uP_64_8853 : std_logic_vector(63 downto 0);
    signal updated_psr_9484 : std_logic_vector(31 downto 0);
    signal updated_y_9559 : std_logic_vector(31 downto 0);
    signal updated_y_9874_delayed_1_0_9772 : std_logic_vector(31 downto 0);
    signal use_alu_add_8605 : std_logic_vector(0 downto 0);
    signal use_alu_add_comp_8709 : std_logic_vector(0 downto 0);
    signal use_alu_and_8605 : std_logic_vector(0 downto 0);
    signal use_alu_div_8605 : std_logic_vector(0 downto 0);
    signal use_alu_mul_8605 : std_logic_vector(0 downto 0);
    signal use_alu_mulscc_8605 : std_logic_vector(0 downto 0);
    signal use_alu_or_8605 : std_logic_vector(0 downto 0);
    signal use_alu_sll_8605 : std_logic_vector(0 downto 0);
    signal use_alu_sra_8605 : std_logic_vector(0 downto 0);
    signal use_alu_srl_8605 : std_logic_vector(0 downto 0);
    signal use_alu_sub_8605 : std_logic_vector(0 downto 0);
    signal use_alu_xnor_8605 : std_logic_vector(0 downto 0);
    signal use_alu_xor_8605 : std_logic_vector(0 downto 0);
    signal uses_iu1_8415 : std_logic_vector(0 downto 0);
    signal valid_bypass_9135 : std_logic_vector(0 downto 0);
    signal wim_8538 : std_logic_vector(31 downto 0);
    signal window_overflow_trap_9618 : std_logic_vector(0 downto 0);
    signal window_underflow_trap_9632 : std_logic_vector(0 downto 0);
    signal with_carry_8605 : std_logic_vector(0 downto 0);
    signal write_asr_8605 : std_logic_vector(0 downto 0);
    signal write_psr_8605 : std_logic_vector(0 downto 0);
    signal write_psr_9570_delayed_1_0_9450 : std_logic_vector(0 downto 0);
    signal write_tbr_8605 : std_logic_vector(0 downto 0);
    signal write_to_psr_8988 : std_logic_vector(0 downto 0);
    signal write_wim_8605 : std_logic_vector(0 downto 0);
    signal write_y_8605 : std_logic_vector(0 downto 0);
    signal y_8544 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    CONCAT_u1_u2_9032_wire_constant <= "00";
    CONCAT_u1_u2_9253_wire_constant <= "00";
    Cmul_8878 <= "0";
    R_ONE_1_8534_wire_constant <= "1";
    R_ZERO_7_9636_wire_constant <= "0000000";
    Vmul_8875 <= "0";
    konst_8368_wire_constant <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000";
    konst_8482_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    konst_8680_wire_constant <= "00000000000000000000000000010111";
    konst_8685_wire_constant <= "00000000000000000000000000010110";
    konst_8690_wire_constant <= "00000000000000000000000000010101";
    konst_8695_wire_constant <= "00000000000000000000000000010100";
    konst_8757_wire_constant <= "00000000000000000000000000000000";
    konst_8763_wire_constant <= "00000000000000000000000000000000";
    konst_8768_wire_constant <= "00000000000000000000000000000000";
    konst_8774_wire_constant <= "00000000000000000000000000000000";
    konst_8782_wire_constant <= "00000000000000000000000000011111";
    konst_8790_wire_constant <= "00000000000000000000000000000000";
    konst_8797_wire_constant <= "0";
    konst_8803_wire_constant <= "0";
    konst_8865_wire_constant <= "00000000000000000000000000011111";
    konst_8870_wire_constant <= "00000000000000000000000000000000";
    konst_8882_wire_constant <= "00000000000000000000000000000000";
    konst_9001_wire_constant <= "00000000000000000000000000000000";
    konst_9005_wire_constant <= "00000000000000000000000000000000";
    konst_9010_wire_constant <= "00000000000000000000000000000000";
    konst_9014_wire_constant <= "00000000000000000000000000000000";
    konst_9199_wire_constant <= "00000000000000000000000000000000";
    konst_9346_wire_constant <= "00000000000000000000000000000000";
    konst_9355_wire_constant <= "00000000000000000000000000000000";
    konst_9359_wire_constant <= "00000000000000000000000000000000";
    konst_9366_wire_constant <= "00000000000000000000000000000000";
    konst_9370_wire_constant <= "00000000000000000000000000000000";
    konst_9375_wire_constant <= "00000000000000000000000000000000";
    konst_9379_wire_constant <= "00000000000000000000000000000000";
    konst_9390_wire_constant <= "00000000000000000000000000000000";
    konst_9491_wire_constant <= "00000000000000000000000000000101";
    konst_9503_wire_constant <= "00000000000000000000000000000101";
    konst_9528_wire_constant <= "00000000000000000000000000000111";
    konst_9548_wire_constant <= "00000000000000000000000000000000";
    konst_9555_wire_constant <= "00000000000000000000000000000000";
    konst_9580_wire_constant <= "00000000000000000000000000000111";
    konst_9624_wire_constant <= "0";
    konst_9628_wire_constant <= "0";
    konst_9848_wire_constant <= "1";
    type_cast_9538_wire_constant <= "01000";
    -- flow-through select operator MUX_8483_inst
    ops_qualified_8484 <= ops_8376 when (get_from_rfile_8647_delayed_1_0_8478(0) /=  '0') else konst_8482_wire_constant;
    -- flow-through select operator MUX_8670_inst
    operand_1_8671 <= pc_8455 when (OR_u1_u1_8667_wire(0) /=  '0') else rf_operand_1_8508;
    -- flow-through select operator MUX_8676_inst
    operand_2_8677 <= imm_operand_8451 when (imm_flag_8403(0) /=  '0') else rf_operand_2_8512;
    -- flow-through select operator MUX_8745_inst
    l_operand_2_8746 <= NOT_u32_u32_8743_wire when (negate_second_operand_8605(0) /=  '0') else operand_2_8677;
    -- flow-through select operator MUX_8758_inst
    MUX_8758_wire <= AND_u32_u32_8756_wire when (use_alu_and_8605(0) /=  '0') else konst_8757_wire_constant;
    -- flow-through select operator MUX_8764_inst
    MUX_8764_wire <= OR_u32_u32_8762_wire when (use_alu_or_8605(0) /=  '0') else konst_8763_wire_constant;
    -- flow-through select operator MUX_8769_inst
    MUX_8769_wire <= i32_xor_result_8751 when (use_alu_xor_8605(0) /=  '0') else konst_8768_wire_constant;
    -- flow-through select operator MUX_8775_inst
    MUX_8775_wire <= XOR_u32_u32_8773_wire when (use_alu_xnor_8605(0) /=  '0') else konst_8774_wire_constant;
    -- flow-through select operator MUX_8785_inst
    Nlogical_8786 <= BITSEL_u32_u1_8783_wire when (issue_logical_8739(0) /=  '0') else Ni_8682;
    -- flow-through select operator MUX_8793_inst
    Zlogical_8794 <= EQ_u32_u1_8791_wire when (issue_logical_8739(0) /=  '0') else Zi_8687;
    -- flow-through select operator MUX_8799_inst
    Vlogical_8800 <= konst_8797_wire_constant when (issue_logical_8739(0) /=  '0') else Vi_8692;
    -- flow-through select operator MUX_8805_inst
    Clogical_8806 <= konst_8803_wire_constant when (issue_logical_8739(0) /=  '0') else Ci_8697;
    -- flow-through select operator MUX_8883_inst
    mul_y_op_1_8884 <= signed_correction_8862 when (signed_mul_div_8605(0) /=  '0') else konst_8882_wire_constant;
    -- flow-through select operator MUX_8995_inst
    MUX_8995_wire <= i32_xor_result_8751 when (write_psr_8605(0) /=  '0') else psr_8516;
    -- flow-through select operator MUX_8996_inst
    post_rett_or_write_psr_psr_8997 <= cti_next_psr_8951 when (exec_rett_8905(0) /=  '0') else MUX_8995_wire;
    -- flow-through select operator MUX_9002_inst
    MUX_9002_wire <= i32_add_sub_result_8727 when (issue_add_sub_8705(0) /=  '0') else konst_9001_wire_constant;
    -- flow-through select operator MUX_9006_inst
    MUX_9006_wire <= i32_logical_op_result_8778 when (issue_logical_8739(0) /=  '0') else konst_9005_wire_constant;
    -- flow-through select operator MUX_9011_inst
    MUX_9011_wire <= imm_operand_8451 when (issue_sethi_8617(0) /=  '0') else konst_9010_wire_constant;
    -- flow-through select operator MUX_9015_inst
    MUX_9015_wire <= i32_shift_result_8823 when (issue_shift_8816(0) /=  '0') else konst_9014_wire_constant;
    -- flow-through select operator MUX_9023_inst
    fast_alu_result_9024 <= i32_mul_result_8857 when (issue_mul_8849(0) /=  '0') else fast_fast_alu_result_9018;
    -- flow-through select operator MUX_9057_inst
    MUX_9057_wire <= CONCAT_u2_u4_9049_wire when (issue_logical_8739(0) /=  '0') else CONCAT_u2_u4_9056_wire;
    -- flow-through select operator MUX_9058_inst
    MUX_9058_wire <= CONCAT_u2_u4_9041_wire when (issue_add_sub_8705(0) /=  '0') else MUX_9057_wire;
    -- flow-through select operator MUX_9059_inst
    fast_alu_cc_flags_9060 <= CONCAT_u2_u4_9033_wire when (issue_mul_8849(0) /=  '0') else MUX_9058_wire;
    -- flow-through select operator MUX_9103_inst
    fast_alu_psr_9104 <= post_rett_or_write_psr_psr_8997 when (write_to_psr_8988(0) /=  '0') else CONCAT_u12_u32_9102_wire;
    -- flow-through select operator MUX_9295_inst
    MUX_9295_wire <= CONCAT_u2_u4_9287_wire when (issue_logical_8739(0) /=  '0') else CONCAT_u2_u4_9294_wire;
    MUX_9296_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_9296_inst_req_0;
      MUX_9296_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_9296_inst_req_1;
      MUX_9296_inst_ack_1<= update_ack(0);
      MUX_9296_inst: SelectSplitProtocol generic map(name => "MUX_9296_inst", data_width => 4, buffering => 1, flow_through => false, full_rate => true) -- 
        port map( x => CONCAT_u2_u4_9279_wire, y => MUX_9295_wire, sel => issue_mulscc_8829, z => MUX_9464_9464_delayed_1_0_9297, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_9312_inst
    MUX_9312_wire <= CONCAT_u2_u4_9310_wire when (issue_div_9432_delayed_1_0_9270(0) /=  '0') else MUX_9464_9464_delayed_1_0_9297;
    -- flow-through select operator MUX_9313_inst
    MUX_9313_wire <= CONCAT_u2_u4_9431_9431_delayed_1_0_9267 when (issue_add_sub_9424_delayed_1_0_9258(0) /=  '0') else MUX_9312_wire;
    -- flow-through select operator MUX_9314_inst
    alu_cc_flags_9315 <= CONCAT_u2_u4_9423_9423_delayed_1_0_9255 when (issue_mul_9416_delayed_1_0_9246(0) /=  '0') else MUX_9313_wire;
    MUX_9347_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_9347_inst_req_0;
      MUX_9347_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_9347_inst_req_1;
      MUX_9347_inst_ack_1<= update_ack(0);
      MUX_9347_inst: SelectSplitProtocol generic map(name => "MUX_9347_inst", data_width => 32, buffering => 1, flow_through => false, full_rate => true) -- 
        port map( x => fast_fast_alu_result_9018, y => konst_9346_wire_constant, sel => OR_u1_u1_9344_wire, z => MUX_9490_9490_delayed_1_0_9348, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_9356_inst
    MUX_9356_wire <= i32_mulscc_result_8843 when (issue_mulscc_8829(0) /=  '0') else konst_9355_wire_constant;
    -- flow-through select operator MUX_9360_inst
    MUX_9360_wire <= psr_8516 when (issue_read_psr_8623(0) /=  '0') else konst_9359_wire_constant;
    -- flow-through select operator MUX_9367_inst
    MUX_9367_wire <= wim_8538 when (issue_read_wim_8629(0) /=  '0') else konst_9366_wire_constant;
    -- flow-through select operator MUX_9371_inst
    MUX_9371_wire <= tbr_8541 when (issue_read_tbr_8635(0) /=  '0') else konst_9370_wire_constant;
    -- flow-through select operator MUX_9376_inst
    MUX_9376_wire <= y_8544 when (issue_read_y_8641(0) /=  '0') else konst_9375_wire_constant;
    -- flow-through select operator MUX_9380_inst
    MUX_9380_wire <= asr_8547 when (issue_read_asr_8647(0) /=  '0') else konst_9379_wire_constant;
    -- flow-through select operator MUX_9391_inst
    MUX_9391_wire <= i32_div_result_9223 when (issue_div_9491_delayed_1_0_9351(0) /=  '0') else konst_9390_wire_constant;
    -- flow-through select operator MUX_9397_inst
    alu_result_9398 <= i32_mul_result_9480_delayed_1_0_9336 when (issue_mul_9479_delayed_1_0_9333(0) /=  '0') else OR_u32_u32_9396_wire;
    -- flow-through select operator MUX_9480_inst
    MUX_9480_wire <= alu_psr_9330 when (OR_u1_u1_9582_9582_delayed_1_0_9466(0) /=  '0') else psr_9584_delayed_1_0_9469;
    -- flow-through select operator MUX_9481_inst
    MUX_9481_wire <= i32_xor_result_9571_delayed_1_0_9453 when (write_psr_9570_delayed_1_0_9450(0) /=  '0') else MUX_9480_wire;
    -- flow-through select operator MUX_9482_inst
    MUX_9482_wire <= cti_next_psr_9569_delayed_1_0_9447 when (exec_rett_9568_delayed_1_0_9444(0) /=  '0') else MUX_9481_wire;
    -- flow-through select operator MUX_9483_inst
    updated_psr_9484 <= psr_9567_delayed_1_0_9441 when (OR_u1_u1_9566_9566_delayed_1_0_9438(0) /=  '0') else MUX_9482_wire;
    -- flow-through select operator MUX_9549_inst
    MUX_9549_wire <= i32_mulscc_y_8843 when (issue_mulscc_8829(0) /=  '0') else konst_9548_wire_constant;
    -- flow-through select operator MUX_9556_inst
    MUX_9556_wire <= i32_xor_result_8751 when (AND_u1_u1_9553_wire(0) /=  '0') else konst_9555_wire_constant;
    -- flow-through select operator MUX_9558_inst
    updated_y_9559 <= i32_mul_y_8893 when (issue_mul_8849(0) /=  '0') else OR_u32_u32_9557_wire;
    -- flow-through select operator MUX_9625_inst
    MUX_9625_wire <= restore_uflow_trap_8555 when (is_restore_8605(0) /=  '0') else konst_9624_wire_constant;
    -- flow-through select operator MUX_9629_inst
    MUX_9629_wire <= cti_window_underflow_trap_8951 when (issue_cti_8929(0) /=  '0') else konst_9628_wire_constant;
    -- flow-through select operator MUX_9637_inst
    ticc_trap_type_9638 <= cti_ticc_trap_type_8951 when (issue_cti_8929(0) /=  '0') else R_ZERO_7_9636_wire_constant;
    -- flow-through slice operator slice_8382_inst
    thread_id_8383 <= exec_info_d_8379(147 downto 144);
    -- flow-through slice operator slice_8386_inst
    stream_id_8387 <= exec_info_d_8379(143 downto 142);
    -- flow-through slice operator slice_8390_inst
    slot_id_8391 <= exec_info_d_8379(141 downto 136);
    -- flow-through slice operator slice_8394_inst
    exec_control_word_8395 <= exec_info_d_8379(135 downto 81);
    -- flow-through slice operator slice_8398_inst
    do_not_bypass_8399 <= exec_info_d_8379(80 downto 80);
    -- flow-through slice operator slice_8402_inst
    imm_flag_8403 <= exec_info_d_8379(79 downto 79);
    -- flow-through slice operator slice_8406_inst
    trap_if_not_super_8407 <= exec_info_d_8379(78 downto 78);
    -- flow-through slice operator slice_8410_inst
    rd_8411 <= exec_info_d_8379(77 downto 73);
    -- flow-through slice operator slice_8414_inst
    uses_iu1_8415 <= exec_info_d_8379(72 downto 72);
    -- flow-through slice operator slice_8418_inst
    send_fast_alu_result_8419 <= exec_info_d_8379(71 downto 71);
    -- flow-through slice operator slice_8422_inst
    iu1_to_iu2_8423 <= exec_info_d_8379(70 downto 70);
    -- flow-through slice operator slice_8426_inst
    iu1_to_sc_8427 <= exec_info_d_8379(69 downto 69);
    -- flow-through slice operator slice_8430_inst
    iu_reg_to_ls_8431 <= exec_info_d_8379(68 downto 68);
    -- flow-through slice operator slice_8434_inst
    iu1_to_ls_trap_8435 <= exec_info_d_8379(67 downto 67);
    -- flow-through slice operator slice_8438_inst
    iu1_to_fu2_8439 <= exec_info_d_8379(66 downto 66);
    -- flow-through slice operator slice_8442_inst
    iu1_to_cu2_8443 <= exec_info_d_8379(65 downto 65);
    -- flow-through slice operator slice_8446_inst
    skip_iu_8447 <= exec_info_d_8379(64 downto 64);
    -- flow-through slice operator slice_8450_inst
    imm_operand_8451 <= exec_info_d_8379(63 downto 32);
    -- flow-through slice operator slice_8454_inst
    pc_8455 <= exec_info_d_8379(31 downto 0);
    -- flow-through slice operator slice_8487_inst
    skip_from_rfile_8488 <= ops_qualified_8484(141 downto 141);
    -- flow-through slice operator slice_8491_inst
    ops_valid_8492 <= ops_qualified_8484(140 downto 140);
    -- flow-through slice operator slice_8495_inst
    thread_id_1_8496 <= ops_qualified_8484(139 downto 136);
    -- flow-through slice operator slice_8499_inst
    stream_id_1_8500 <= ops_qualified_8484(135 downto 134);
    -- flow-through slice operator slice_8503_inst
    slot_id_1_8504 <= ops_qualified_8484(133 downto 128);
    -- flow-through slice operator slice_8507_inst
    rf_operand_1_8508 <= ops_qualified_8484(127 downto 96);
    -- flow-through slice operator slice_8511_inst
    rf_operand_2_8512 <= ops_qualified_8484(95 downto 64);
    -- flow-through slice operator slice_8515_inst
    psr_8516 <= ops_qualified_8484(63 downto 32);
    -- flow-through slice operator slice_8519_inst
    sreg_value_8520 <= ops_qualified_8484(31 downto 0);
    -- flow-through slice operator slice_8856_inst
    i32_mul_result_8857 <= uP_64_8853(31 downto 0);
    -- flow-through slice operator slice_8887_inst
    mul_y_op_2_8888 <= uP_64_8853(63 downto 32);
    -- flow-through slice operator slice_9097_inst
    slice_9097_wire <= psr_8516(31 downto 24);
    -- flow-through slice operator slice_9101_inst
    slice_9101_wire <= psr_8516(19 downto 0);
    slice_9318_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_9318_inst_req_0;
      slice_9318_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_9318_inst_req_1;
      slice_9318_inst_ack_1<= update_ack(0);
      slice_9318_inst: SliceSplitProtocol generic map(name => "slice_9318_inst", in_data_width => 32, high_index => 31, low_index => 24, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => psr_8516, dout => slice_9471_9471_delayed_1_0_9319, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_9322_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_9322_inst_req_0;
      slice_9322_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_9322_inst_req_1;
      slice_9322_inst_ack_1<= update_ack(0);
      slice_9322_inst: SliceSplitProtocol generic map(name => "slice_9322_inst", in_data_width => 32, high_index => 19, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => psr_8516, dout => slice_9475_9475_delayed_1_0_9323, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through slice operator slice_9516_inst
    iu_proc_ilvl_9517 <= post_rett_or_write_psr_psr_8997(11 downto 8);
    -- flow-through slice operator slice_9536_inst
    slice_9536_wire <= post_rett_or_write_psr_psr_8997(4 downto 0);
    -- interlock W_asr_8545_inst
    process(sreg_value_8520) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sreg_value_8520(31 downto 0);
      asr_8547 <= tmp_var; -- 
    end process;
    W_cti_next_psr_9569_delayed_1_0_9445_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_cti_next_psr_9569_delayed_1_0_9445_inst_req_0;
      W_cti_next_psr_9569_delayed_1_0_9445_inst_ack_0<= wack(0);
      rreq(0) <= W_cti_next_psr_9569_delayed_1_0_9445_inst_req_1;
      W_cti_next_psr_9569_delayed_1_0_9445_inst_ack_1<= rack(0);
      W_cti_next_psr_9569_delayed_1_0_9445_inst : InterlockBuffer generic map ( -- 
        name => "W_cti_next_psr_9569_delayed_1_0_9445_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cti_next_psr_8951,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => cti_next_psr_9569_delayed_1_0_9447,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_exec_info_d_8377_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_exec_info_d_8377_inst_req_0;
      W_exec_info_d_8377_inst_ack_0<= wack(0);
      rreq(0) <= W_exec_info_d_8377_inst_req_1;
      W_exec_info_d_8377_inst_ack_1<= rack(0);
      W_exec_info_d_8377_inst : InterlockBuffer generic map ( -- 
        name => "W_exec_info_d_8377_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 150,
        out_data_width => 150,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => exec_info_8365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => exec_info_d_8379,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_exec_rett_9568_delayed_1_0_9442_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_exec_rett_9568_delayed_1_0_9442_inst_req_0;
      W_exec_rett_9568_delayed_1_0_9442_inst_ack_0<= wack(0);
      rreq(0) <= W_exec_rett_9568_delayed_1_0_9442_inst_req_1;
      W_exec_rett_9568_delayed_1_0_9442_inst_ack_1<= rack(0);
      W_exec_rett_9568_delayed_1_0_9442_inst : InterlockBuffer generic map ( -- 
        name => "W_exec_rett_9568_delayed_1_0_9442_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => exec_rett_8905,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => exec_rett_9568_delayed_1_0_9444,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_get_from_rfile_8647_delayed_1_0_8476_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_get_from_rfile_8647_delayed_1_0_8476_inst_req_0;
      W_get_from_rfile_8647_delayed_1_0_8476_inst_ack_0<= wack(0);
      rreq(0) <= W_get_from_rfile_8647_delayed_1_0_8476_inst_req_1;
      W_get_from_rfile_8647_delayed_1_0_8476_inst_ack_1<= rack(0);
      W_get_from_rfile_8647_delayed_1_0_8476_inst : InterlockBuffer generic map ( -- 
        name => "W_get_from_rfile_8647_delayed_1_0_8476_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => get_from_rfile_8370,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => get_from_rfile_8647_delayed_1_0_8478,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_i32_mul_result_9480_delayed_1_0_9334_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_i32_mul_result_9480_delayed_1_0_9334_inst_req_0;
      W_i32_mul_result_9480_delayed_1_0_9334_inst_ack_0<= wack(0);
      rreq(0) <= W_i32_mul_result_9480_delayed_1_0_9334_inst_req_1;
      W_i32_mul_result_9480_delayed_1_0_9334_inst_ack_1<= rack(0);
      W_i32_mul_result_9480_delayed_1_0_9334_inst : InterlockBuffer generic map ( -- 
        name => "W_i32_mul_result_9480_delayed_1_0_9334_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i32_mul_result_8857,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => i32_mul_result_9480_delayed_1_0_9336,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_i32_xor_result_9571_delayed_1_0_9451_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_i32_xor_result_9571_delayed_1_0_9451_inst_req_0;
      W_i32_xor_result_9571_delayed_1_0_9451_inst_ack_0<= wack(0);
      rreq(0) <= W_i32_xor_result_9571_delayed_1_0_9451_inst_req_1;
      W_i32_xor_result_9571_delayed_1_0_9451_inst_ack_1<= rack(0);
      W_i32_xor_result_9571_delayed_1_0_9451_inst : InterlockBuffer generic map ( -- 
        name => "W_i32_xor_result_9571_delayed_1_0_9451_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i32_xor_result_8751,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => i32_xor_result_9571_delayed_1_0_9453,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_issue_add_sub_9424_delayed_1_0_9256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_issue_add_sub_9424_delayed_1_0_9256_inst_req_0;
      W_issue_add_sub_9424_delayed_1_0_9256_inst_ack_0<= wack(0);
      rreq(0) <= W_issue_add_sub_9424_delayed_1_0_9256_inst_req_1;
      W_issue_add_sub_9424_delayed_1_0_9256_inst_ack_1<= rack(0);
      W_issue_add_sub_9424_delayed_1_0_9256_inst : InterlockBuffer generic map ( -- 
        name => "W_issue_add_sub_9424_delayed_1_0_9256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => issue_add_sub_8705,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => issue_add_sub_9424_delayed_1_0_9258,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_issue_div_9432_delayed_1_0_9268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_issue_div_9432_delayed_1_0_9268_inst_req_0;
      W_issue_div_9432_delayed_1_0_9268_inst_ack_0<= wack(0);
      rreq(0) <= W_issue_div_9432_delayed_1_0_9268_inst_req_1;
      W_issue_div_9432_delayed_1_0_9268_inst_ack_1<= rack(0);
      W_issue_div_9432_delayed_1_0_9268_inst : InterlockBuffer generic map ( -- 
        name => "W_issue_div_9432_delayed_1_0_9268_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => issue_div_9211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => issue_div_9432_delayed_1_0_9270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_issue_div_9491_delayed_1_0_9349_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_issue_div_9491_delayed_1_0_9349_inst_req_0;
      W_issue_div_9491_delayed_1_0_9349_inst_ack_0<= wack(0);
      rreq(0) <= W_issue_div_9491_delayed_1_0_9349_inst_req_1;
      W_issue_div_9491_delayed_1_0_9349_inst_ack_1<= rack(0);
      W_issue_div_9491_delayed_1_0_9349_inst : InterlockBuffer generic map ( -- 
        name => "W_issue_div_9491_delayed_1_0_9349_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => issue_div_9211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => issue_div_9491_delayed_1_0_9351,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_issue_mul_9416_delayed_1_0_9244_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_issue_mul_9416_delayed_1_0_9244_inst_req_0;
      W_issue_mul_9416_delayed_1_0_9244_inst_ack_0<= wack(0);
      rreq(0) <= W_issue_mul_9416_delayed_1_0_9244_inst_req_1;
      W_issue_mul_9416_delayed_1_0_9244_inst_ack_1<= rack(0);
      W_issue_mul_9416_delayed_1_0_9244_inst : InterlockBuffer generic map ( -- 
        name => "W_issue_mul_9416_delayed_1_0_9244_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => issue_mul_8849,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => issue_mul_9416_delayed_1_0_9246,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_issue_mul_9479_delayed_1_0_9331_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_issue_mul_9479_delayed_1_0_9331_inst_req_0;
      W_issue_mul_9479_delayed_1_0_9331_inst_ack_0<= wack(0);
      rreq(0) <= W_issue_mul_9479_delayed_1_0_9331_inst_req_1;
      W_issue_mul_9479_delayed_1_0_9331_inst_ack_1<= rack(0);
      W_issue_mul_9479_delayed_1_0_9331_inst : InterlockBuffer generic map ( -- 
        name => "W_issue_mul_9479_delayed_1_0_9331_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => issue_mul_8849,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => issue_mul_9479_delayed_1_0_9333,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_iu_to_fu_trapped_9827_inst
    process(trap_or_error_9816) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := trap_or_error_9816(0 downto 0);
      iu_to_fu_trapped_9829 <= tmp_var; -- 
    end process;
    -- interlock W_iu_to_ls_trapped_9817_inst
    process(trap_or_error_9816) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := trap_or_error_9816(0 downto 0);
      iu_to_ls_trapped_9819 <= tmp_var; -- 
    end process;
    W_psr_9567_delayed_1_0_9439_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_psr_9567_delayed_1_0_9439_inst_req_0;
      W_psr_9567_delayed_1_0_9439_inst_ack_0<= wack(0);
      rreq(0) <= W_psr_9567_delayed_1_0_9439_inst_req_1;
      W_psr_9567_delayed_1_0_9439_inst_ack_1<= rack(0);
      W_psr_9567_delayed_1_0_9439_inst : InterlockBuffer generic map ( -- 
        name => "W_psr_9567_delayed_1_0_9439_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => psr_8516,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => psr_9567_delayed_1_0_9441,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_psr_9584_delayed_1_0_9467_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_psr_9584_delayed_1_0_9467_inst_req_0;
      W_psr_9584_delayed_1_0_9467_inst_ack_0<= wack(0);
      rreq(0) <= W_psr_9584_delayed_1_0_9467_inst_req_1;
      W_psr_9584_delayed_1_0_9467_inst_ack_1<= rack(0);
      W_psr_9584_delayed_1_0_9467_inst : InterlockBuffer generic map ( -- 
        name => "W_psr_9584_delayed_1_0_9467_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => psr_8516,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => psr_9584_delayed_1_0_9469,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_send_to_sc_9697_inst
    process(iu1_to_sc_8427) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := iu1_to_sc_8427(0 downto 0);
      send_to_sc_9699 <= tmp_var; -- 
    end process;
    -- interlock W_send_to_wb_9751_inst
    process(iu1_to_iu2_8423) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := iu1_to_iu2_8423(0 downto 0);
      send_to_wb_9753 <= tmp_var; -- 
    end process;
    W_send_to_wb_9880_delayed_1_0_9784_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send_to_wb_9880_delayed_1_0_9784_inst_req_0;
      W_send_to_wb_9880_delayed_1_0_9784_inst_ack_0<= wack(0);
      rreq(0) <= W_send_to_wb_9880_delayed_1_0_9784_inst_req_1;
      W_send_to_wb_9880_delayed_1_0_9784_inst_ack_1<= rack(0);
      W_send_to_wb_9880_delayed_1_0_9784_inst : InterlockBuffer generic map ( -- 
        name => "W_send_to_wb_9880_delayed_1_0_9784_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send_to_wb_9753,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send_to_wb_9880_delayed_1_0_9786,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_tbr_8539_inst
    process(sreg_value_8520) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sreg_value_8520(31 downto 0);
      tbr_8541 <= tmp_var; -- 
    end process;
    W_updated_y_9874_delayed_1_0_9770_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_updated_y_9874_delayed_1_0_9770_inst_req_0;
      W_updated_y_9874_delayed_1_0_9770_inst_ack_0<= wack(0);
      rreq(0) <= W_updated_y_9874_delayed_1_0_9770_inst_req_1;
      W_updated_y_9874_delayed_1_0_9770_inst_ack_1<= rack(0);
      W_updated_y_9874_delayed_1_0_9770_inst : InterlockBuffer generic map ( -- 
        name => "W_updated_y_9874_delayed_1_0_9770_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => updated_y_9559,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => updated_y_9874_delayed_1_0_9772,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_wim_8536_inst
    process(sreg_value_8520) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sreg_value_8520(31 downto 0);
      wim_8538 <= tmp_var; -- 
    end process;
    W_write_psr_9570_delayed_1_0_9448_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_psr_9570_delayed_1_0_9448_inst_req_0;
      W_write_psr_9570_delayed_1_0_9448_inst_ack_0<= wack(0);
      rreq(0) <= W_write_psr_9570_delayed_1_0_9448_inst_req_1;
      W_write_psr_9570_delayed_1_0_9448_inst_ack_1<= rack(0);
      W_write_psr_9570_delayed_1_0_9448_inst : InterlockBuffer generic map ( -- 
        name => "W_write_psr_9570_delayed_1_0_9448_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_psr_8605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_psr_9570_delayed_1_0_9450,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_y_8542_inst
    process(sreg_value_8520) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sreg_value_8520(31 downto 0);
      y_8544 <= tmp_var; -- 
    end process;
    do_while_stmt_8361_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_9848_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_8361_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_8361_branch_req_0,
          ack0 => do_while_stmt_8361_branch_ack_0,
          ack1 => do_while_stmt_8361_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator ADD_u32_u32_8892_inst
    i32_mul_y_8893 <= std_logic_vector(unsigned(mul_y_op_1_8884) + unsigned(mul_y_op_2_8888));
    -- flow through binary operator AND_u1_u1_8616_inst
    issue_sethi_8617 <= (NOT_u1_u1_8614_wire and is_sethi_8605);
    -- flow through binary operator AND_u1_u1_8622_inst
    issue_read_psr_8623 <= (NOT_u1_u1_8620_wire and read_psr_8605);
    -- flow through binary operator AND_u1_u1_8628_inst
    issue_read_wim_8629 <= (NOT_u1_u1_8626_wire and read_wim_8605);
    -- flow through binary operator AND_u1_u1_8634_inst
    issue_read_tbr_8635 <= (NOT_u1_u1_8632_wire and read_tbr_8605);
    -- flow through binary operator AND_u1_u1_8640_inst
    issue_read_y_8641 <= (NOT_u1_u1_8638_wire and read_y_8605);
    -- flow through binary operator AND_u1_u1_8646_inst
    issue_read_asr_8647 <= (NOT_u1_u1_8644_wire and read_asr_8605);
    -- flow through binary operator AND_u1_u1_8704_inst
    issue_add_sub_8705 <= (NOT_u1_u1_8700_wire and OR_u1_u1_8703_wire);
    -- flow through binary operator AND_u1_u1_8738_inst
    issue_logical_8739 <= (NOT_u1_u1_8730_wire and OR_u1_u1_8737_wire);
    -- flow through binary operator AND_u1_u1_8815_inst
    issue_shift_8816 <= (NOT_u1_u1_8809_wire and OR_u1_u1_8814_wire);
    -- flow through binary operator AND_u1_u1_8828_inst
    issue_mulscc_8829 <= (NOT_u1_u1_8826_wire and use_alu_mulscc_8605);
    -- flow through binary operator AND_u1_u1_8848_inst
    issue_mul_8849 <= (NOT_u1_u1_8846_wire and use_alu_mul_8605);
    -- flow through binary operator AND_u1_u1_8898_inst
    exec_call_8899 <= (NOT_u1_u1_8896_wire and is_call_8605);
    -- flow through binary operator AND_u1_u1_8904_inst
    exec_rett_8905 <= (NOT_u1_u1_8902_wire and is_rett_8605);
    -- flow through binary operator AND_u1_u1_8910_inst
    exec_jmpl_8911 <= (NOT_u1_u1_8908_wire and is_jmpl_8605);
    -- flow through binary operator AND_u1_u1_8916_inst
    exec_ticc_8917 <= (NOT_u1_u1_8914_wire and is_ticc_8605);
    -- flow through binary operator AND_u1_u1_8922_inst
    exec_bicc_8923 <= (NOT_u1_u1_8920_wire and is_bicc_8605);
    -- flow through binary operator AND_u1_u1_8928_inst
    issue_cti_8929 <= (NOT_u1_u1_8926_wire and cti_8605);
    -- flow through binary operator AND_u1_u1_8955_inst
    cti_trap_8956 <= (issue_cti_8929 and cti_trap_status_8951);
    -- flow through binary operator AND_u1_u1_8987_inst
    write_to_psr_8988 <= (NOT_u1_u1_8983_wire and OR_u1_u1_8986_wire);
    -- flow through binary operator AND_u1_u1_9066_inst
    AND_u1_u1_9066_wire <= (NOT_u1_u1_9063_wire and NOT_u1_u1_9065_wire);
    -- flow through binary operator AND_u1_u1_9073_inst
    AND_u1_u1_9073_wire <= (OR_u1_u1_9071_wire and set_cc_8605);
    -- flow through binary operator AND_u1_u1_9076_inst
    fast_update_psr_9077 <= (AND_u1_u1_9066_wire and OR_u1_u1_9075_wire);
    -- flow through binary operator AND_u1_u1_9083_inst
    AND_u1_u1_9083_wire <= (NOT_u1_u1_9080_wire and NOT_u1_u1_9082_wire);
    -- flow through binary operator AND_u1_u1_9090_inst
    AND_u1_u1_9090_wire <= (set_cc_8605 and OR_u1_u1_9089_wire);
    -- flow through binary operator AND_u1_u1_9091_inst
    send_cc_bypass_9092 <= (AND_u1_u1_9083_wire and AND_u1_u1_9090_wire);
    -- flow through binary operator AND_u1_u1_9110_inst
    AND_u1_u1_9110_wire <= (NOT_u1_u1_9107_wire and NOT_u1_u1_9109_wire);
    -- flow through binary operator AND_u1_u1_9112_inst
    send_alu_bypass_9113 <= (AND_u1_u1_9110_wire and send_fast_alu_result_8419);
    -- flow through binary operator AND_u1_u1_9197_inst
    AND_u1_u1_9197_wire <= (NOT_u1_u1_9195_wire and use_alu_div_8605);
    -- flow through binary operator AND_u1_u1_9201_inst
    div_by_0_trap_9202 <= (AND_u1_u1_9197_wire and EQ_u32_u1_9200_wire);
    -- flow through binary operator AND_u1_u1_9207_inst
    AND_u1_u1_9207_wire <= (NOT_u1_u1_9205_wire and use_alu_div_8605);
    -- flow through binary operator AND_u1_u1_9210_inst
    issue_div_9211 <= (AND_u1_u1_9207_wire and NOT_u1_u1_9209_wire);
    -- flow through binary operator AND_u1_u1_9240_inst
    AND_u1_u1_9240_wire <= (issue_add_sub_8705 and i32_add_sub_ovflow_trap_8727);
    -- flow through binary operator AND_u1_u1_9464_inst
    AND_u1_u1_9464_wire <= (set_cc_8605 and OR_u1_u1_9463_wire);
    -- flow through binary operator AND_u1_u1_9493_inst
    AND_u1_u1_9493_wire <= (write_psr_8605 and BITSEL_u32_u1_9492_wire);
    -- flow through binary operator AND_u1_u1_9495_inst
    iu_enable_traps_9496 <= (NOT_u1_u1_9487_wire and OR_u1_u1_9494_wire);
    -- flow through binary operator AND_u1_u1_9501_inst
    AND_u1_u1_9501_wire <= (NOT_u1_u1_9499_wire and write_psr_8605);
    -- flow through binary operator AND_u1_u1_9506_inst
    iu_disable_traps_9507 <= (AND_u1_u1_9501_wire and NOT_u1_u1_9505_wire);
    -- flow through binary operator AND_u1_u1_9512_inst
    iu_set_proc_ilvl_9513 <= (NOT_u1_u1_9510_wire and write_psr_8605);
    -- flow through binary operator AND_u1_u1_9524_inst
    iu_set_S_9525 <= (NOT_u1_u1_9520_wire and OR_u1_u1_9523_wire);
    -- flow through binary operator AND_u1_u1_9540_inst
    AND_u1_u1_9540_wire <= (write_to_psr_8988 and UGE_u5_u1_9539_wire);
    -- flow through binary operator AND_u1_u1_9541_inst
    sr_illegal_instr_trap_9542 <= (NOT_u1_u1_9533_wire and AND_u1_u1_9540_wire);
    -- flow through binary operator AND_u1_u1_9553_inst
    AND_u1_u1_9553_wire <= (NOT_u1_u1_9551_wire and write_y_8605);
    -- flow through binary operator AND_u1_u1_9566_inst
    AND_u1_u1_9566_wire <= (issue_cti_8929 and cti_illegal_instr_trap_8951);
    -- flow through binary operator AND_u1_u1_9568_inst
    illegal_instr_trap_9569 <= (NOT_u1_u1_9562_wire and OR_u1_u1_9567_wire);
    -- flow through binary operator AND_u1_u1_9589_inst
    AND_u1_u1_9589_wire <= (trap_if_not_super_8407 and NOT_u1_u1_9588_wire);
    -- flow through binary operator AND_u1_u1_9592_inst
    AND_u1_u1_9592_wire <= (issue_cti_8929 and cti_privileged_instr_trap_8951);
    -- flow through binary operator AND_u1_u1_9594_inst
    priv_instr_trap_9595 <= (NOT_u1_u1_9585_wire and OR_u1_u1_9593_wire);
    -- flow through binary operator AND_u1_u1_9599_inst
    alu_overflow_trap_9600 <= (issue_add_sub_8705 and i32_add_sub_ovflow_trap_8727);
    -- flow through binary operator AND_u1_u1_9604_inst
    trap_instr_trap_9605 <= (issue_cti_8929 and cti_trap_instr_trap_8951);
    -- flow through binary operator AND_u1_u1_9609_inst
    mem_addr_not_aligned_trap_9610 <= (issue_cti_8929 and cti_mem_address_not_aligned_trap_8951);
    -- flow through binary operator AND_u1_u1_9616_inst
    AND_u1_u1_9616_wire <= (is_save_8605 and save_ovflow_trap_8551);
    -- flow through binary operator AND_u1_u1_9617_inst
    window_overflow_trap_9618 <= (NOT_u1_u1_9613_wire and AND_u1_u1_9616_wire);
    -- flow through binary operator AND_u1_u1_9631_inst
    window_underflow_trap_9632 <= (NOT_u1_u1_9621_wire and OR_u1_u1_9630_wire);
    -- flow through binary operator AND_u1_u1_9680_inst
    AND_u1_u1_9680_wire <= (issue_cti_8929 and cti_processor_error_mode_8951);
    -- flow through binary operator AND_u1_u1_9685_inst
    exec_processor_error_mode_9686 <= (NOT_u1_u1_9677_wire and OR_u1_u1_9684_wire);
    -- flow through binary operator AND_u1_u1_9690_inst
    br_taken_9691 <= (issue_cti_8929 and cti_br_taken_8951);
    -- flow through binary operator AND_u1_u1_9695_inst
    annul_next_9696 <= (issue_cti_8929 and cti_annul_next_8951);
    -- flow through binary operator AND_u32_u32_8756_inst
    AND_u32_u32_8756_wire <= (operand_1_8671 and l_operand_2_8746);
    -- flow through binary operator BITSEL_u150_u1_8369_inst
    process(exec_info_8365) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(exec_info_8365, konst_8368_wire_constant, tmp_var);
      get_from_rfile_8370 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_8681_inst
    process(psr_8516) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(psr_8516, konst_8680_wire_constant, tmp_var);
      Ni_8682 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_8686_inst
    process(psr_8516) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(psr_8516, konst_8685_wire_constant, tmp_var);
      Zi_8687 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_8691_inst
    process(psr_8516) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(psr_8516, konst_8690_wire_constant, tmp_var);
      Vi_8692 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_8696_inst
    process(psr_8516) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(psr_8516, konst_8695_wire_constant, tmp_var);
      Ci_8697 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_8783_inst
    process(i32_logical_op_result_8778) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(i32_logical_op_result_8778, konst_8782_wire_constant, tmp_var);
      BITSEL_u32_u1_8783_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_8866_inst
    process(i32_mul_result_8857) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(i32_mul_result_8857, konst_8865_wire_constant, tmp_var);
      Nmul_8867 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_9492_inst
    process(post_rett_or_write_psr_psr_8997) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(post_rett_or_write_psr_psr_8997, konst_9491_wire_constant, tmp_var);
      BITSEL_u32_u1_9492_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_9504_inst
    process(post_rett_or_write_psr_psr_8997) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(post_rett_or_write_psr_psr_8997, konst_9503_wire_constant, tmp_var);
      BITSEL_u32_u1_9504_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_9529_inst
    process(post_rett_or_write_psr_psr_8997) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(post_rett_or_write_psr_psr_8997, konst_9528_wire_constant, tmp_var);
      iu_S_9530 <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_9581_inst
    process(psr_8516) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(psr_8516, konst_9580_wire_constant, tmp_var);
      S_9582 <= tmp_var; --
    end process;
    -- shared split operator group (70) : CONCAT_u12_u14_9763_inst 
    ApConcat_group_70: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u6_u12_9759_wire & CONCAT_u1_u2_9762_wire;
      CONCAT_u12_u14_9868_9868_delayed_1_0_9764 <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u12_u14_9763_inst_req_0;
      CONCAT_u12_u14_9763_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u12_u14_9763_inst_req_1;
      CONCAT_u12_u14_9763_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_70_gI: SplitGuardInterface generic map(name => "ApConcat_group_70_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_70",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 2, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- flow through binary operator CONCAT_u12_u32_9102_inst
    process(CONCAT_u8_u12_9099_wire, slice_9101_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u12_9099_wire, slice_9101_wire, tmp_var);
      CONCAT_u12_u32_9102_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u12_u32_9329_inst
    process(CONCAT_u8_u12_9327_wire, slice_9475_9475_delayed_1_0_9323) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u12_9327_wire, slice_9475_9475_delayed_1_0_9323, tmp_var);
      alu_psr_9330 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u13_u109_9179_inst
    process(CONCAT_u6_u13_9173_wire, CONCAT_u64_u96_9178_wire) -- 
      variable tmp_var : std_logic_vector(108 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u6_u13_9173_wire, CONCAT_u64_u96_9178_wire, tmp_var);
      fast_result_to_wb_9180 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u13_u20_9715_inst
    process(CONCAT_u6_u13_9707_wire, CONCAT_u2_u7_9714_wire) -- 
      variable tmp_var : std_logic_vector(19 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u6_u13_9707_wire, CONCAT_u2_u7_9714_wire, tmp_var);
      CONCAT_u13_u20_9715_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u13_u83_9129_inst
    process(CONCAT_u5_u13_9121_wire, CONCAT_u6_u70_9128_wire) -- 
      variable tmp_var : std_logic_vector(82 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u5_u13_9121_wire, CONCAT_u6_u70_9128_wire, tmp_var);
      bypass_to_reg_file_9130 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u14_u126_9782_inst
    process(CONCAT_u12_u14_9868_9868_delayed_1_0_9764, CONCAT_u48_u112_9781_wire) -- 
      variable tmp_var : std_logic_vector(125 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u12_u14_9868_9868_delayed_1_0_9764, CONCAT_u48_u112_9781_wire, tmp_var);
      to_iu_wb_9783 <= tmp_var; --
    end process;
    -- shared split operator group (77) : CONCAT_u15_u16_9768_inst 
    ApConcat_group_77: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= traps_9657 & skip_iu_8447;
      CONCAT_u15_u16_9871_9871_delayed_1_0_9769 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u15_u16_9768_inst_req_0;
      CONCAT_u15_u16_9768_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u15_u16_9768_inst_req_1;
      CONCAT_u15_u16_9768_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_77_gI: SplitGuardInterface generic map(name => "ApConcat_group_77_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_77",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 77
    -- flow through binary operator CONCAT_u16_u48_9777_inst
    process(CONCAT_u15_u16_9871_9871_delayed_1_0_9769, updated_psr_9484) -- 
      variable tmp_var : std_logic_vector(47 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u15_u16_9871_9871_delayed_1_0_9769, updated_psr_9484, tmp_var);
      CONCAT_u16_u48_9777_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9029_inst
    process(Nmul_8867, Zmul_8872) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Nmul_8867, Zmul_8872, tmp_var);
      CONCAT_u1_u2_9029_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9037_inst
    process(Naddsub_8727, Zaddsub_8727) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Naddsub_8727, Zaddsub_8727, tmp_var);
      CONCAT_u1_u2_9037_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9040_inst
    process(Vaddsub_8727, Caddsub_8727) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Vaddsub_8727, Caddsub_8727, tmp_var);
      CONCAT_u1_u2_9040_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9045_inst
    process(Nlogical_8786, Zlogical_8794) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Nlogical_8786, Zlogical_8794, tmp_var);
      CONCAT_u1_u2_9045_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9048_inst
    process(Vlogical_8800, Clogical_8806) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Vlogical_8800, Clogical_8806, tmp_var);
      CONCAT_u1_u2_9048_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9052_inst
    process(Ni_8682, Zi_8687) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Ni_8682, Zi_8687, tmp_var);
      CONCAT_u1_u2_9052_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9055_inst
    process(Vi_8692, Ci_8697) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Vi_8692, Ci_8697, tmp_var);
      CONCAT_u1_u2_9055_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9250_inst
    process(Nmul_8867, Zmul_8872) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Nmul_8867, Zmul_8872, tmp_var);
      CONCAT_u1_u2_9250_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9262_inst
    process(Naddsub_8727, Zaddsub_8727) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Naddsub_8727, Zaddsub_8727, tmp_var);
      CONCAT_u1_u2_9262_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9265_inst
    process(Vaddsub_8727, Caddsub_8727) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Vaddsub_8727, Caddsub_8727, tmp_var);
      CONCAT_u1_u2_9265_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9275_inst
    process(Nmulscc_8843, Zmulscc_8843) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Nmulscc_8843, Zmulscc_8843, tmp_var);
      CONCAT_u1_u2_9275_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9278_inst
    process(Vmulscc_8843, Cmulscc_8843) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Vmulscc_8843, Cmulscc_8843, tmp_var);
      CONCAT_u1_u2_9278_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9283_inst
    process(Nlogical_8786, Zlogical_8794) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Nlogical_8786, Zlogical_8794, tmp_var);
      CONCAT_u1_u2_9283_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9286_inst
    process(Vlogical_8800, Clogical_8806) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Vlogical_8800, Clogical_8806, tmp_var);
      CONCAT_u1_u2_9286_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9290_inst
    process(Ni_8682, Zi_8687) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Ni_8682, Zi_8687, tmp_var);
      CONCAT_u1_u2_9290_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9293_inst
    process(Vi_8692, Ci_8697) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Vi_8692, Ci_8697, tmp_var);
      CONCAT_u1_u2_9293_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9306_inst
    process(Ndiv_9223, Zdiv_9223) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Ndiv_9223, Zdiv_9223, tmp_var);
      CONCAT_u1_u2_9306_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9309_inst
    process(Vdiv_9223, Cdiv_9223) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(Vdiv_9223, Cdiv_9223, tmp_var);
      CONCAT_u1_u2_9309_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9642_inst
    process(illegal_instr_trap_9569, priv_instr_trap_9595) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(illegal_instr_trap_9569, priv_instr_trap_9595, tmp_var);
      CONCAT_u1_u2_9642_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9647_inst
    process(div_by_0_trap_9202, trap_instr_trap_9605) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(div_by_0_trap_9202, trap_instr_trap_9605, tmp_var);
      CONCAT_u1_u2_9647_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9651_inst
    process(mem_addr_not_aligned_trap_9610, window_underflow_trap_9632) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(mem_addr_not_aligned_trap_9610, window_underflow_trap_9632, tmp_var);
      CONCAT_u1_u2_9651_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9710_inst
    process(iu_enable_traps_9496, iu_disable_traps_9507) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(iu_enable_traps_9496, iu_disable_traps_9507, tmp_var);
      CONCAT_u1_u2_9710_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9718_inst
    process(iu_set_S_9525, iu_S_9530) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(iu_set_S_9525, iu_S_9530, tmp_var);
      CONCAT_u1_u2_9718_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9721_inst
    process(br_taken_9691, annul_next_9696) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(br_taken_9691, annul_next_9696, tmp_var);
      CONCAT_u1_u2_9721_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9725_inst
    process(exec_processor_error_mode_9686, iunit_has_trapped_9674) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(exec_processor_error_mode_9686, iunit_has_trapped_9674, tmp_var);
      CONCAT_u1_u2_9725_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_9762_inst
    process(exec_processor_error_mode_9686, iunit_has_trapped_9674) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(exec_processor_error_mode_9686, iunit_has_trapped_9674, tmp_var);
      CONCAT_u1_u2_9762_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u5_9117_inst
    process(send_alu_bypass_9113, thread_id_8383) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApConcat_proc(send_alu_bypass_9113, thread_id_8383, tmp_var);
      CONCAT_u1_u5_9117_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u5_9149_inst
    process(send_cc_bypass_9092, thread_id_8383) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApConcat_proc(send_cc_bypass_9092, thread_id_8383, tmp_var);
      CONCAT_u1_u5_9149_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u5_9713_inst
    process(iu_set_proc_ilvl_9513, iu_proc_ilvl_9517) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApConcat_proc(iu_set_proc_ilvl_9513, iu_proc_ilvl_9517, tmp_var);
      CONCAT_u1_u5_9713_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u6_9124_inst
    process(fast_update_psr_9077, rd_8411) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(fast_update_psr_9077, rd_8411, tmp_var);
      CONCAT_u1_u6_9124_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u8_9654_inst
    process(window_overflow_trap_9618, ticc_trap_type_9638) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(window_overflow_trap_9618, ticc_trap_type_9638, tmp_var);
      CONCAT_u1_u8_9654_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u20_u90_9731_inst
    process(CONCAT_u13_u20_9715_wire, CONCAT_u4_u70_9730_wire) -- 
      variable tmp_var : std_logic_vector(89 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u13_u20_9715_wire, CONCAT_u4_u70_9730_wire, tmp_var);
      to_sc_9732 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u10_9655_inst
    process(CONCAT_u1_u2_9651_wire, CONCAT_u1_u8_9654_wire) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9651_wire, CONCAT_u1_u8_9654_wire, tmp_var);
      CONCAT_u2_u10_9655_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u3_9644_inst
    process(CONCAT_u1_u2_9642_wire, alu_overflow_trap_9600) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9642_wire, alu_overflow_trap_9600, tmp_var);
      CONCAT_u2_u3_9644_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u4_9033_inst
    process(CONCAT_u1_u2_9029_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9029_wire, CONCAT_u1_u2_9032_wire_constant, tmp_var);
      CONCAT_u2_u4_9033_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u4_9041_inst
    process(CONCAT_u1_u2_9037_wire, CONCAT_u1_u2_9040_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9037_wire, CONCAT_u1_u2_9040_wire, tmp_var);
      CONCAT_u2_u4_9041_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u4_9049_inst
    process(CONCAT_u1_u2_9045_wire, CONCAT_u1_u2_9048_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9045_wire, CONCAT_u1_u2_9048_wire, tmp_var);
      CONCAT_u2_u4_9049_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u4_9056_inst
    process(CONCAT_u1_u2_9052_wire, CONCAT_u1_u2_9055_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9052_wire, CONCAT_u1_u2_9055_wire, tmp_var);
      CONCAT_u2_u4_9056_wire <= tmp_var; --
    end process;
    -- shared split operator group (117) : CONCAT_u2_u4_9254_inst 
    ApConcat_group_117: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u2_9250_wire;
      CONCAT_u2_u4_9423_9423_delayed_1_0_9255 <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u2_u4_9254_inst_req_0;
      CONCAT_u2_u4_9254_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u2_u4_9254_inst_req_1;
      CONCAT_u2_u4_9254_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_117_gI: SplitGuardInterface generic map(name => "ApConcat_group_117_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_117",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "00",
          constant_width => 2,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 117
    -- shared split operator group (118) : CONCAT_u2_u4_9266_inst 
    ApConcat_group_118: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u2_9262_wire & CONCAT_u1_u2_9265_wire;
      CONCAT_u2_u4_9431_9431_delayed_1_0_9267 <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u2_u4_9266_inst_req_0;
      CONCAT_u2_u4_9266_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u2_u4_9266_inst_req_1;
      CONCAT_u2_u4_9266_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_118_gI: SplitGuardInterface generic map(name => "ApConcat_group_118_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_118",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 2, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 118
    -- flow through binary operator CONCAT_u2_u4_9279_inst
    process(CONCAT_u1_u2_9275_wire, CONCAT_u1_u2_9278_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9275_wire, CONCAT_u1_u2_9278_wire, tmp_var);
      CONCAT_u2_u4_9279_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u4_9287_inst
    process(CONCAT_u1_u2_9283_wire, CONCAT_u1_u2_9286_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9283_wire, CONCAT_u1_u2_9286_wire, tmp_var);
      CONCAT_u2_u4_9287_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u4_9294_inst
    process(CONCAT_u1_u2_9290_wire, CONCAT_u1_u2_9293_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9290_wire, CONCAT_u1_u2_9293_wire, tmp_var);
      CONCAT_u2_u4_9294_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u4_9310_inst
    process(CONCAT_u1_u2_9306_wire, CONCAT_u1_u2_9309_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9306_wire, CONCAT_u1_u2_9309_wire, tmp_var);
      CONCAT_u2_u4_9310_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u4_9722_inst
    process(CONCAT_u1_u2_9718_wire, CONCAT_u1_u2_9721_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9718_wire, CONCAT_u1_u2_9721_wire, tmp_var);
      CONCAT_u2_u4_9722_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u66_9729_inst
    process(CONCAT_u1_u2_9725_wire, CONCAT_u32_u64_9728_wire) -- 
      variable tmp_var : std_logic_vector(65 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9725_wire, CONCAT_u32_u64_9728_wire, tmp_var);
      CONCAT_u2_u66_9729_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u7_9714_inst
    process(CONCAT_u1_u2_9710_wire, CONCAT_u1_u5_9713_wire) -- 
      variable tmp_var : std_logic_vector(6 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9710_wire, CONCAT_u1_u5_9713_wire, tmp_var);
      CONCAT_u2_u7_9714_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u2_u8_9120_inst
    process(stream_id_8387, slot_id_8391) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(stream_id_8387, slot_id_8391, tmp_var);
      CONCAT_u2_u8_9120_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u32_u64_9127_inst
    process(fast_alu_psr_9104, fast_alu_result_9024) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(fast_alu_psr_9104, fast_alu_result_9024, tmp_var);
      CONCAT_u32_u64_9127_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u32_u64_9176_inst
    process(fast_alu_psr_9104, fast_alu_result_9024) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(fast_alu_psr_9104, fast_alu_result_9024, tmp_var);
      CONCAT_u32_u64_9176_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u32_u64_9728_inst
    process(i32_add_sub_result_8727, post_rett_or_write_psr_psr_8997) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(i32_add_sub_result_8727, post_rett_or_write_psr_psr_8997, tmp_var);
      CONCAT_u32_u64_9728_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u32_u64_9780_inst
    process(updated_y_9874_delayed_1_0_9772, alu_result_9398) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(updated_y_9874_delayed_1_0_9772, alu_result_9398, tmp_var);
      CONCAT_u32_u64_9780_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u3_u5_9648_inst
    process(CONCAT_u2_u3_9644_wire, CONCAT_u1_u2_9647_wire) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u3_9644_wire, CONCAT_u1_u2_9647_wire, tmp_var);
      CONCAT_u3_u5_9648_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u48_u112_9781_inst
    process(CONCAT_u16_u48_9777_wire, CONCAT_u32_u64_9780_wire) -- 
      variable tmp_var : std_logic_vector(111 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u16_u48_9777_wire, CONCAT_u32_u64_9780_wire, tmp_var);
      CONCAT_u48_u112_9781_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u4_u6_9169_inst
    process(thread_id_8383, stream_id_8387) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(thread_id_8383, stream_id_8387, tmp_var);
      CONCAT_u4_u6_9169_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u4_u6_9703_inst
    process(thread_id_8383, stream_id_8387) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(thread_id_8383, stream_id_8387, tmp_var);
      CONCAT_u4_u6_9703_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u4_u6_9757_inst
    process(thread_id_8383, stream_id_8387) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(thread_id_8383, stream_id_8387, tmp_var);
      CONCAT_u4_u6_9757_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u4_u6_9833_inst
    process(thread_id_8383, stream_id_8387) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(thread_id_8383, stream_id_8387, tmp_var);
      CONCAT_u4_u6_9833_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u4_u70_9730_inst
    process(CONCAT_u2_u4_9722_wire, CONCAT_u2_u66_9729_wire) -- 
      variable tmp_var : std_logic_vector(69 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u4_9722_wire, CONCAT_u2_u66_9729_wire, tmp_var);
      CONCAT_u4_u70_9730_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u5_u13_9121_inst
    process(CONCAT_u1_u5_9117_wire, CONCAT_u2_u8_9120_wire) -- 
      variable tmp_var : std_logic_vector(12 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u5_9117_wire, CONCAT_u2_u8_9120_wire, tmp_var);
      CONCAT_u5_u13_9121_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u5_u15_9656_inst
    process(CONCAT_u3_u5_9648_wire, CONCAT_u2_u10_9655_wire) -- 
      variable tmp_var : std_logic_vector(14 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u3_u5_9648_wire, CONCAT_u2_u10_9655_wire, tmp_var);
      traps_9657 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u5_u7_9151_inst
    process(CONCAT_u1_u5_9149_wire, stream_id_8387) -- 
      variable tmp_var : std_logic_vector(6 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u5_9149_wire, stream_id_8387, tmp_var);
      CONCAT_u5_u7_9151_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u64_u96_9178_inst
    process(CONCAT_u32_u64_9176_wire, i32_mul_y_8893) -- 
      variable tmp_var : std_logic_vector(95 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u32_u64_9176_wire, i32_mul_y_8893, tmp_var);
      CONCAT_u64_u96_9178_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u6_u10_9154_inst
    process(slot_id_8391, fast_alu_cc_flags_9060) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApConcat_proc(slot_id_8391, fast_alu_cc_flags_9060, tmp_var);
      CONCAT_u6_u10_9154_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u6_u12_9759_inst
    process(CONCAT_u4_u6_9757_wire, slot_id_8391) -- 
      variable tmp_var : std_logic_vector(11 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u4_u6_9757_wire, slot_id_8391, tmp_var);
      CONCAT_u6_u12_9759_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u6_u13_9173_inst
    process(CONCAT_u4_u6_9169_wire, CONCAT_u6_u7_9172_wire) -- 
      variable tmp_var : std_logic_vector(12 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u4_u6_9169_wire, CONCAT_u6_u7_9172_wire, tmp_var);
      CONCAT_u6_u13_9173_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u6_u13_9707_inst
    process(CONCAT_u4_u6_9703_wire, CONCAT_u6_u7_9706_wire) -- 
      variable tmp_var : std_logic_vector(12 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u4_u6_9703_wire, CONCAT_u6_u7_9706_wire, tmp_var);
      CONCAT_u6_u13_9707_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u6_u13_9837_inst
    process(CONCAT_u4_u6_9833_wire, CONCAT_u6_u7_9836_wire) -- 
      variable tmp_var : std_logic_vector(12 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u4_u6_9833_wire, CONCAT_u6_u7_9836_wire, tmp_var);
      to_fpu_9838 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u6_u70_9128_inst
    process(CONCAT_u1_u6_9124_wire, CONCAT_u32_u64_9127_wire) -- 
      variable tmp_var : std_logic_vector(69 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u6_9124_wire, CONCAT_u32_u64_9127_wire, tmp_var);
      CONCAT_u6_u70_9128_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u6_u7_9172_inst
    process(slot_id_8391, fast_update_psr_9077) -- 
      variable tmp_var : std_logic_vector(6 downto 0); -- 
    begin -- 
      ApConcat_proc(slot_id_8391, fast_update_psr_9077, tmp_var);
      CONCAT_u6_u7_9172_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u6_u7_9706_inst
    process(slot_id_8391, skip_iu_8447) -- 
      variable tmp_var : std_logic_vector(6 downto 0); -- 
    begin -- 
      ApConcat_proc(slot_id_8391, skip_iu_8447, tmp_var);
      CONCAT_u6_u7_9706_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u6_u7_9836_inst
    process(slot_id_8391, iu_to_fu_trapped_9829) -- 
      variable tmp_var : std_logic_vector(6 downto 0); -- 
    begin -- 
      ApConcat_proc(slot_id_8391, iu_to_fu_trapped_9829, tmp_var);
      CONCAT_u6_u7_9836_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u7_u17_9155_inst
    process(CONCAT_u5_u7_9151_wire, CONCAT_u6_u10_9154_wire) -- 
      variable tmp_var : std_logic_vector(16 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u5_u7_9151_wire, CONCAT_u6_u10_9154_wire, tmp_var);
      bypass_cc_to_reg_file_9156 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u8_u12_9099_inst
    process(slice_9097_wire, fast_alu_cc_flags_9060) -- 
      variable tmp_var : std_logic_vector(11 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_9097_wire, fast_alu_cc_flags_9060, tmp_var);
      CONCAT_u8_u12_9099_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u8_u12_9327_inst
    process(slice_9471_9471_delayed_1_0_9319, alu_cc_flags_9315) -- 
      variable tmp_var : std_logic_vector(11 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_9471_9471_delayed_1_0_9319, alu_cc_flags_9315, tmp_var);
      CONCAT_u8_u12_9327_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_8791_inst
    process(i32_logical_op_result_8778) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(i32_logical_op_result_8778, konst_8790_wire_constant, tmp_var);
      EQ_u32_u1_8791_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_8871_inst
    process(i32_mul_result_8857) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(i32_mul_result_8857, konst_8870_wire_constant, tmp_var);
      Zmul_8872 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_9200_inst
    process(operand_2_8677) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(operand_2_8677, konst_9199_wire_constant, tmp_var);
      EQ_u32_u1_9200_wire <= tmp_var; --
    end process;
    -- flow through binary operator NEQ_u6_u1_9683_inst
    process(slot_id_8391, slot_id_1_8504) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(slot_id_8391, slot_id_1_8504, tmp_var);
      NEQ_u6_u1_9683_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_8609_inst
    process(uses_iu1_8415) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", uses_iu1_8415, tmp_var);
      NOT_u1_u1_8609_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8614_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8614_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8620_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8620_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8626_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8626_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8632_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8632_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8638_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8638_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8644_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8644_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8700_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8700_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8708_inst
    process(use_alu_add_8605) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", use_alu_add_8605, tmp_var);
      use_alu_add_comp_8709 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8730_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8730_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8809_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8809_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8826_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8826_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8846_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8846_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8896_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8896_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8902_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8902_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8908_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8908_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8914_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8914_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8920_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8920_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8926_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8926_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_8983_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_8983_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9063_inst
    process(skip_iu_8447) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_iu_8447, tmp_var);
      NOT_u1_u1_9063_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9065_inst
    process(do_not_bypass_8399) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", do_not_bypass_8399, tmp_var);
      NOT_u1_u1_9065_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9080_inst
    process(skip_iu_8447) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_iu_8447, tmp_var);
      NOT_u1_u1_9080_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9082_inst
    process(do_not_bypass_8399) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", do_not_bypass_8399, tmp_var);
      NOT_u1_u1_9082_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9107_inst
    process(skip_iu_8447) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_iu_8447, tmp_var);
      NOT_u1_u1_9107_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9109_inst
    process(do_not_bypass_8399) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", do_not_bypass_8399, tmp_var);
      NOT_u1_u1_9109_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9195_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_9195_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9205_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_9205_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9209_inst
    process(div_by_0_trap_9202) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", div_by_0_trap_9202, tmp_var);
      NOT_u1_u1_9209_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9487_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_9487_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9499_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_9499_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9505_inst
    process(BITSEL_u32_u1_9504_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_9504_wire, tmp_var);
      NOT_u1_u1_9505_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9510_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_9510_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9520_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_9520_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9533_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_9533_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9551_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_9551_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9562_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_9562_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9585_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_9585_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9588_inst
    process(S_9582) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", S_9582, tmp_var);
      NOT_u1_u1_9588_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9613_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_9613_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9621_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_9621_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_9677_inst
    process(skip_alu_exec_8611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_alu_exec_8611, tmp_var);
      NOT_u1_u1_9677_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u32_u32_8743_inst
    process(operand_2_8677) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", operand_2_8677, tmp_var);
      NOT_u32_u32_8743_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_8610_inst
    skip_alu_exec_8611 <= (skip_iu_8447 or NOT_u1_u1_8609_wire);
    -- flow through binary operator OR_u1_u1_8663_inst
    OR_u1_u1_8663_wire <= (is_call_8605 or is_bicc_8605);
    -- flow through binary operator OR_u1_u1_8666_inst
    OR_u1_u1_8666_wire <= (is_fbfcc_8605 or is_cbccc_8605);
    -- flow through binary operator OR_u1_u1_8667_inst
    OR_u1_u1_8667_wire <= (OR_u1_u1_8663_wire or OR_u1_u1_8666_wire);
    -- flow through binary operator OR_u1_u1_8703_inst
    OR_u1_u1_8703_wire <= (use_alu_sub_8605 or use_alu_add_8605);
    -- flow through binary operator OR_u1_u1_8733_inst
    OR_u1_u1_8733_wire <= (use_alu_and_8605 or use_alu_or_8605);
    -- flow through binary operator OR_u1_u1_8736_inst
    OR_u1_u1_8736_wire <= (use_alu_xor_8605 or use_alu_xnor_8605);
    -- flow through binary operator OR_u1_u1_8737_inst
    OR_u1_u1_8737_wire <= (OR_u1_u1_8733_wire or OR_u1_u1_8736_wire);
    -- flow through binary operator OR_u1_u1_8812_inst
    OR_u1_u1_8812_wire <= (use_alu_sll_8605 or use_alu_srl_8605);
    -- flow through binary operator OR_u1_u1_8814_inst
    OR_u1_u1_8814_wire <= (OR_u1_u1_8812_wire or use_alu_sra_8605);
    -- flow through binary operator OR_u1_u1_8986_inst
    OR_u1_u1_8986_wire <= (write_psr_8605 or exec_rett_8905);
    -- flow through binary operator OR_u1_u1_9069_inst
    OR_u1_u1_9069_wire <= (issue_add_sub_8705 or issue_logical_8739);
    -- flow through binary operator OR_u1_u1_9071_inst
    OR_u1_u1_9071_wire <= (OR_u1_u1_9069_wire or issue_mul_8849);
    -- flow through binary operator OR_u1_u1_9075_inst
    OR_u1_u1_9075_wire <= (AND_u1_u1_9073_wire or write_to_psr_8988);
    -- flow through binary operator OR_u1_u1_9087_inst
    OR_u1_u1_9087_wire <= (issue_add_sub_8705 or issue_logical_8739);
    -- flow through binary operator OR_u1_u1_9089_inst
    OR_u1_u1_9089_wire <= (OR_u1_u1_9087_wire or issue_mul_8849);
    -- flow through binary operator OR_u1_u1_9134_inst
    valid_bypass_9135 <= (send_alu_bypass_9113 or fast_update_psr_9077);
    -- flow through binary operator OR_u1_u1_9227_inst
    OR_u1_u1_9227_wire <= (issue_add_sub_8705 or issue_mul_8849);
    -- flow through binary operator OR_u1_u1_9229_inst
    OR_u1_u1_9229_wire <= (OR_u1_u1_9227_wire or issue_div_9211);
    -- flow through binary operator OR_u1_u1_9232_inst
    OR_u1_u1_9232_wire <= (issue_mulscc_8829 or issue_logical_8739);
    -- flow through binary operator OR_u1_u1_9234_inst
    OR_u1_u1_9234_wire <= (OR_u1_u1_9232_wire or issue_shift_8816);
    -- flow through binary operator OR_u1_u1_9235_inst
    alu_was_used_9236 <= (OR_u1_u1_9229_wire or OR_u1_u1_9234_wire);
    -- flow through binary operator OR_u1_u1_9242_inst
    alu_trap_9243 <= (AND_u1_u1_9240_wire or div_by_0_trap_9202);
    -- flow through binary operator OR_u1_u1_9340_inst
    OR_u1_u1_9340_wire <= (issue_add_sub_8705 or issue_shift_8816);
    -- flow through binary operator OR_u1_u1_9343_inst
    OR_u1_u1_9343_wire <= (issue_logical_8739 or issue_sethi_8617);
    -- flow through binary operator OR_u1_u1_9344_inst
    OR_u1_u1_9344_wire <= (OR_u1_u1_9340_wire or OR_u1_u1_9343_wire);
    -- shared split operator group (227) : OR_u1_u1_9437_inst 
    ApIntOr_group_227: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= alu_trap_9243 & cti_trap_8956;
      OR_u1_u1_9566_9566_delayed_1_0_9438 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u1_u1_9437_inst_req_0;
      OR_u1_u1_9437_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u1_u1_9437_inst_req_1;
      OR_u1_u1_9437_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_227_gI: SplitGuardInterface generic map(name => "ApIntOr_group_227_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_227",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 227
    -- flow through binary operator OR_u1_u1_9459_inst
    OR_u1_u1_9459_wire <= (issue_add_sub_8705 or issue_div_9211);
    -- flow through binary operator OR_u1_u1_9462_inst
    OR_u1_u1_9462_wire <= (issue_mul_8849 or issue_logical_8739);
    -- flow through binary operator OR_u1_u1_9463_inst
    OR_u1_u1_9463_wire <= (OR_u1_u1_9459_wire or OR_u1_u1_9462_wire);
    -- shared split operator group (231) : OR_u1_u1_9465_inst 
    ApIntOr_group_231: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= issue_mulscc_8829 & AND_u1_u1_9464_wire;
      OR_u1_u1_9582_9582_delayed_1_0_9466 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u1_u1_9465_inst_req_0;
      OR_u1_u1_9465_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u1_u1_9465_inst_req_1;
      OR_u1_u1_9465_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_231_gI: SplitGuardInterface generic map(name => "ApIntOr_group_231_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_231",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 231
    -- flow through binary operator OR_u1_u1_9494_inst
    OR_u1_u1_9494_wire <= (exec_rett_8905 or AND_u1_u1_9493_wire);
    -- flow through binary operator OR_u1_u1_9523_inst
    OR_u1_u1_9523_wire <= (write_psr_8605 or exec_rett_8905);
    -- flow through binary operator OR_u1_u1_9567_inst
    OR_u1_u1_9567_wire <= (sr_illegal_instr_trap_9542 or AND_u1_u1_9566_wire);
    -- flow through binary operator OR_u1_u1_9593_inst
    OR_u1_u1_9593_wire <= (AND_u1_u1_9589_wire or AND_u1_u1_9592_wire);
    -- flow through binary operator OR_u1_u1_9630_inst
    OR_u1_u1_9630_wire <= (MUX_9625_wire or MUX_9629_wire);
    -- flow through binary operator OR_u1_u1_9661_inst
    OR_u1_u1_9661_wire <= (illegal_instr_trap_9569 or priv_instr_trap_9595);
    -- flow through binary operator OR_u1_u1_9664_inst
    OR_u1_u1_9664_wire <= (alu_overflow_trap_9600 or div_by_0_trap_9202);
    -- flow through binary operator OR_u1_u1_9665_inst
    OR_u1_u1_9665_wire <= (OR_u1_u1_9661_wire or OR_u1_u1_9664_wire);
    -- flow through binary operator OR_u1_u1_9668_inst
    OR_u1_u1_9668_wire <= (trap_instr_trap_9605 or mem_addr_not_aligned_trap_9610);
    -- flow through binary operator OR_u1_u1_9671_inst
    OR_u1_u1_9671_wire <= (window_underflow_trap_9632 or window_overflow_trap_9618);
    -- flow through binary operator OR_u1_u1_9672_inst
    OR_u1_u1_9672_wire <= (OR_u1_u1_9668_wire or OR_u1_u1_9671_wire);
    -- flow through binary operator OR_u1_u1_9673_inst
    iunit_has_trapped_9674 <= (OR_u1_u1_9665_wire or OR_u1_u1_9672_wire);
    -- flow through binary operator OR_u1_u1_9684_inst
    OR_u1_u1_9684_wire <= (AND_u1_u1_9680_wire or NEQ_u6_u1_9683_wire);
    -- flow through binary operator OR_u1_u1_9815_inst
    trap_or_error_9816 <= (iunit_has_trapped_9674 or exec_processor_error_mode_9686);
    -- flow through binary operator OR_u32_u32_8762_inst
    OR_u32_u32_8762_wire <= (operand_1_8671 or l_operand_2_8746);
    -- flow through binary operator OR_u32_u32_8765_inst
    OR_u32_u32_8765_wire <= (MUX_8758_wire or MUX_8764_wire);
    -- flow through binary operator OR_u32_u32_8776_inst
    OR_u32_u32_8776_wire <= (MUX_8769_wire or MUX_8775_wire);
    -- flow through binary operator OR_u32_u32_8777_inst
    i32_logical_op_result_8778 <= (OR_u32_u32_8765_wire or OR_u32_u32_8776_wire);
    -- flow through binary operator OR_u32_u32_9007_inst
    OR_u32_u32_9007_wire <= (MUX_9002_wire or MUX_9006_wire);
    -- flow through binary operator OR_u32_u32_9016_inst
    OR_u32_u32_9016_wire <= (MUX_9011_wire or MUX_9015_wire);
    -- flow through binary operator OR_u32_u32_9017_inst
    fast_fast_alu_result_9018 <= (OR_u32_u32_9007_wire or OR_u32_u32_9016_wire);
    -- shared split operator group (253) : OR_u32_u32_9361_inst 
    ApIntOr_group_253: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= MUX_9356_wire & MUX_9360_wire;
      OR_u32_u32_9504_9504_delayed_1_0_9362 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_9361_inst_req_0;
      OR_u32_u32_9361_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_9361_inst_req_1;
      OR_u32_u32_9361_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_253_gI: SplitGuardInterface generic map(name => "ApIntOr_group_253_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_253",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 253
    -- flow through binary operator OR_u32_u32_9372_inst
    OR_u32_u32_9372_wire <= (MUX_9367_wire or MUX_9371_wire);
    -- flow through binary operator OR_u32_u32_9381_inst
    OR_u32_u32_9381_wire <= (MUX_9376_wire or MUX_9380_wire);
    -- shared split operator group (256) : OR_u32_u32_9382_inst 
    ApIntOr_group_256: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= OR_u32_u32_9372_wire & OR_u32_u32_9381_wire;
      OR_u32_u32_9524_9524_delayed_1_0_9383 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_9382_inst_req_0;
      OR_u32_u32_9382_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_9382_inst_req_1;
      OR_u32_u32_9382_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_256_gI: SplitGuardInterface generic map(name => "ApIntOr_group_256_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_256",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 256
    -- flow through binary operator OR_u32_u32_9392_inst
    OR_u32_u32_9392_wire <= (MUX_9490_9490_delayed_1_0_9348 or MUX_9391_wire);
    -- flow through binary operator OR_u32_u32_9394_inst
    OR_u32_u32_9394_wire <= (OR_u32_u32_9392_wire or OR_u32_u32_9504_9504_delayed_1_0_9362);
    -- flow through binary operator OR_u32_u32_9396_inst
    OR_u32_u32_9396_wire <= (OR_u32_u32_9394_wire or OR_u32_u32_9524_9524_delayed_1_0_9383);
    -- flow through binary operator OR_u32_u32_9557_inst
    OR_u32_u32_9557_wire <= (MUX_9549_wire or MUX_9556_wire);
    -- flow through binary operator UGE_u5_u1_9539_inst
    process(slice_9536_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(slice_9536_wire, type_cast_9538_wire_constant, tmp_var);
      UGE_u5_u1_9539_wire <= tmp_var; --
    end process;
    -- flow through binary operator XOR_u32_u32_8750_inst
    i32_xor_result_8751 <= (operand_1_8671 xor l_operand_2_8746);
    -- flow through binary operator XOR_u32_u32_8773_inst
    XOR_u32_u32_8773_wire <= not (operand_1_8671 xor l_operand_2_8746);
    -- shared inport operator group (0) : RPIPE_iunit_register_file_read_access_response_8375_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(141 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_iunit_register_file_read_access_response_8375_inst_req_0;
      RPIPE_iunit_register_file_read_access_response_8375_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_iunit_register_file_read_access_response_8375_inst_req_1;
      RPIPE_iunit_register_file_read_access_response_8375_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= get_from_rfile_8370(0);
      ops_8376 <= data_out(141 downto 0);
      iunit_register_file_read_access_response_read_0_gI: SplitGuardInterface generic map(name => "iunit_register_file_read_access_response_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      iunit_register_file_read_access_response_read_0: InputPort_P2P -- 
        generic map ( name => "iunit_register_file_read_access_response_read_0", data_width => 142,    bypass_flag => false,   	nonblocking_read_flag => false,  barrier_flag => false,   queue_depth =>  2)
        port map (-- 
          sample_req => reqL(0) , 
          sample_ack => ackL(0), 
          update_req => reqR(0), 
          update_ack => ackR(0), 
          data => data_out, 
          oreq => iunit_register_file_read_access_response_pipe_read_req(0),
          oack => iunit_register_file_read_access_response_pipe_read_ack(0),
          odata => iunit_register_file_read_access_response_pipe_read_data(141 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_teu_idispatch_to_iunit_exec_8364_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(149 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_teu_idispatch_to_iunit_exec_8364_inst_req_0;
      RPIPE_teu_idispatch_to_iunit_exec_8364_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_teu_idispatch_to_iunit_exec_8364_inst_req_1;
      RPIPE_teu_idispatch_to_iunit_exec_8364_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      exec_info_8365 <= data_out(149 downto 0);
      teu_idispatch_to_iunit_exec_read_1_gI: SplitGuardInterface generic map(name => "teu_idispatch_to_iunit_exec_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      teu_idispatch_to_iunit_exec_read_1: InputPort_P2P -- 
        generic map ( name => "teu_idispatch_to_iunit_exec_read_1", data_width => 150,    bypass_flag => false,   	nonblocking_read_flag => false,  barrier_flag => false,   queue_depth =>  2)
        port map (-- 
          sample_req => reqL(0) , 
          sample_ack => ackL(0), 
          update_req => reqR(0), 
          update_ack => ackR(0), 
          data => data_out, 
          oreq => teu_idispatch_to_iunit_exec_pipe_read_req(0),
          oack => teu_idispatch_to_iunit_exec_pipe_read_ack(0),
          odata => teu_idispatch_to_iunit_exec_pipe_read_data(149 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(108 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_inst_req_0;
      WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_inst_req_1;
      WPIPE_iunit_exec_fast_alu_result_to_writeback_9182_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_fast_alu_result_8419(0);
      data_in <= fast_result_to_wb_9180;
      iunit_exec_fast_alu_result_to_writeback_write_0_gI: SplitGuardInterface generic map(name => "iunit_exec_fast_alu_result_to_writeback_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      iunit_exec_fast_alu_result_to_writeback_write_0: OutputPortRevised -- 
        generic map ( name => "iunit_exec_fast_alu_result_to_writeback", data_width => 109, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => iunit_exec_fast_alu_result_to_writeback_pipe_write_req(0),
          oack => iunit_exec_fast_alu_result_to_writeback_pipe_write_ack(0),
          odata => iunit_exec_fast_alu_result_to_writeback_pipe_write_data(108 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_iunit_exec_to_writeback_9788_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(125 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_iunit_exec_to_writeback_9788_inst_req_0;
      WPIPE_iunit_exec_to_writeback_9788_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_iunit_exec_to_writeback_9788_inst_req_1;
      WPIPE_iunit_exec_to_writeback_9788_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_wb_9880_delayed_1_0_9786(0);
      data_in <= to_iu_wb_9783;
      iunit_exec_to_writeback_write_1_gI: SplitGuardInterface generic map(name => "iunit_exec_to_writeback_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      iunit_exec_to_writeback_write_1: OutputPortRevised -- 
        generic map ( name => "iunit_exec_to_writeback", data_width => 126, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => iunit_exec_to_writeback_pipe_write_req(0),
          oack => iunit_exec_to_writeback_pipe_write_ack(0),
          odata => iunit_exec_to_writeback_pipe_write_data(125 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(16 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_inst_req_0;
      WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_inst_req_1;
      WPIPE_noblock_iunit_exec_bypass_cc_signal_to_register_file_9157_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= bypass_cc_to_reg_file_9156;
      noblock_iunit_exec_bypass_cc_signal_to_register_file_write_2_gI: SplitGuardInterface generic map(name => "noblock_iunit_exec_bypass_cc_signal_to_register_file_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_iunit_exec_bypass_cc_signal_to_register_file_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_iunit_exec_bypass_cc_signal_to_register_file", data_width => 17, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_req(0),
          oack => noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_ack(0),
          odata => noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_data(16 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(82 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_inst_req_0;
      WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_inst_req_1;
      WPIPE_noblock_iunit_exec_bypass_signal_to_register_file_9136_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= bypass_to_reg_file_9130;
      noblock_iunit_exec_bypass_signal_to_register_file_write_3_gI: SplitGuardInterface generic map(name => "noblock_iunit_exec_bypass_signal_to_register_file_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_iunit_exec_bypass_signal_to_register_file_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_iunit_exec_bypass_signal_to_register_file", data_width => 83, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_req(0),
          oack => noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_ack(0),
          odata => noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_data(82 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_inst_req_0;
      WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_inst_req_1;
      WPIPE_noblock_iunit_exec_to_regfile_credit_return_8533_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= ops_valid_8492(0);
      data_in <= R_ONE_1_8534_wire_constant;
      noblock_iunit_exec_to_regfile_credit_return_write_4_gI: SplitGuardInterface generic map(name => "noblock_iunit_exec_to_regfile_credit_return_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_iunit_exec_to_regfile_credit_return_write_4: OutputPortRevised -- 
        generic map ( name => "noblock_iunit_exec_to_regfile_credit_return", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_iunit_exec_to_regfile_credit_return_pipe_write_req(0),
          oack => noblock_iunit_exec_to_regfile_credit_return_pipe_write_ack(0),
          odata => noblock_iunit_exec_to_regfile_credit_return_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_teu_iunit_to_stream_corrector_9734_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(89 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_teu_iunit_to_stream_corrector_9734_inst_req_0;
      WPIPE_teu_iunit_to_stream_corrector_9734_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_teu_iunit_to_stream_corrector_9734_inst_req_1;
      WPIPE_teu_iunit_to_stream_corrector_9734_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_sc_9699(0);
      data_in <= to_sc_9732;
      teu_iunit_to_stream_corrector_write_5_gI: SplitGuardInterface generic map(name => "teu_iunit_to_stream_corrector_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      teu_iunit_to_stream_corrector_write_5: OutputPortRevised -- 
        generic map ( name => "teu_iunit_to_stream_corrector", data_width => 90, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => teu_iunit_to_stream_corrector_pipe_write_req(0),
          oack => teu_iunit_to_stream_corrector_pipe_write_ack(0),
          odata => teu_iunit_to_stream_corrector_pipe_write_data(89 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared outport operator group (6) : WPIPE_teu_iunit_trap_to_fpunit_9840_inst 
    OutportGroup_6: Block -- 
      signal data_in: std_logic_vector(12 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_teu_iunit_trap_to_fpunit_9840_inst_req_0;
      WPIPE_teu_iunit_trap_to_fpunit_9840_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_teu_iunit_trap_to_fpunit_9840_inst_req_1;
      WPIPE_teu_iunit_trap_to_fpunit_9840_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= iu1_to_fu2_8439(0);
      data_in <= to_fpu_9838;
      teu_iunit_trap_to_fpunit_write_6_gI: SplitGuardInterface generic map(name => "teu_iunit_trap_to_fpunit_write_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      teu_iunit_trap_to_fpunit_write_6: OutputPortRevised -- 
        generic map ( name => "teu_iunit_trap_to_fpunit", data_width => 13, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => teu_iunit_trap_to_fpunit_pipe_write_req(0),
          oack => teu_iunit_trap_to_fpunit_pipe_write_ack(0),
          odata => teu_iunit_trap_to_fpunit_pipe_write_data(12 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 6
    -- shared outport operator group (7) : WPIPE_teu_iunit_trap_to_loadstore_9821_inst 
    OutportGroup_7: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_teu_iunit_trap_to_loadstore_9821_inst_req_0;
      WPIPE_teu_iunit_trap_to_loadstore_9821_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_teu_iunit_trap_to_loadstore_9821_inst_req_1;
      WPIPE_teu_iunit_trap_to_loadstore_9821_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= iu1_to_ls_trap_8435(0);
      data_in <= iu_to_ls_trapped_9819;
      teu_iunit_trap_to_loadstore_write_7_gI: SplitGuardInterface generic map(name => "teu_iunit_trap_to_loadstore_write_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      teu_iunit_trap_to_loadstore_write_7: OutputPortRevised -- 
        generic map ( name => "teu_iunit_trap_to_loadstore", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => teu_iunit_trap_to_loadstore_pipe_write_req(0),
          oack => teu_iunit_trap_to_loadstore_pipe_write_ack(0),
          odata => teu_iunit_trap_to_loadstore_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 7
    volatile_operator_save_window_trap_8862: save_window_trap_Volatile port map(psr => psr_8516, wim => wim_8538, ovflow_trap => save_ovflow_trap_8551); 
    volatile_operator_restore_window_trap_8863: restore_window_trap_Volatile port map(psr => psr_8516, wim => wim_8538, uflow_trap => restore_uflow_trap_8555); 
    volatile_operator_decode_alu_exec_control_word_8864: decode_alu_exec_control_word_Volatile port map(cw => exec_control_word_8395, cti => cti_8605, is_call => is_call_8605, is_jmpl => is_jmpl_8605, is_rett => is_rett_8605, is_bicc => is_bicc_8605, is_fbfcc => is_fbfcc_8605, is_cbccc => is_cbccc_8605, is_ticc => is_ticc_8605, annul_flag => annul_flag_8605, br_cond => br_cond_8605, alu => alu_8605, use_alu_add => use_alu_add_8605, is_alu_sub => use_alu_sub_8605, is_alu_mul => use_alu_mul_8605, is_alu_mulscc => use_alu_mulscc_8605, is_alu_div => use_alu_div_8605, is_alu_sll => use_alu_sll_8605, is_alu_srl => use_alu_srl_8605, is_alu_sra => use_alu_sra_8605, is_alu_and => use_alu_and_8605, is_alu_or => use_alu_or_8605, use_alu_xor => use_alu_xor_8605, is_alu_xnor => use_alu_xnor_8605, signed_mul_div => signed_mul_div_8605, negate_second_operand => negate_second_operand_8605, with_carry => with_carry_8605, set_cc => set_cc_8605, tagged_alu_op => tagged_alu_op_8605, trap_on_overflow => trap_on_overflow_8605, misc => misc_8605, is_sethi => is_sethi_8605, write_psr => write_psr_8605, write_wim => write_wim_8605, write_tbr => write_tbr_8605, write_y => write_y_8605, write_asr => write_asr_8605, read_psr => read_psr_8605, read_wim => read_wim_8605, read_tbr => read_tbr_8605, read_y => read_y_8605, read_asr => read_asr_8605, asr_id => asr_id_8605, is_save => is_save_8605, is_restore => is_restore_8605, dti => dti_8605, is_iu_dti => iu_dti_8605, is_load_to_debug => is_load_to_debug_8605, is_store_to_debug => is_store_to_debug_8605); 
    volatile_operator_i32_add_sub_8892: i32_add_sub_Volatile port map(subtract_flag => use_alu_add_comp_8709, with_carry => with_carry_8605, set_cc => set_cc_8605, tagged_op => tagged_alu_op_8605, trap_on_ovflow => trap_on_overflow_8605, Ni => Ni_8682, Zi => Zi_8687, Vi => Vi_8692, Ci => Ci_8697, x => operand_1_8671, y => operand_2_8677, result => i32_add_sub_result_8727, No => Naddsub_8727, Zo => Zaddsub_8727, Vo => Vaddsub_8727, Co => Caddsub_8727, overflow_trap => i32_add_sub_ovflow_trap_8727); 
    volatile_operator_i32_shift_8921: i32_shift_Volatile port map(is_sll => use_alu_sll_8605, is_srl => use_alu_srl_8605, is_sra => use_alu_sra_8605, x => operand_1_8671, shift_amount => operand_2_8677, result => i32_shift_result_8823); 
    volatile_operator_i32_mulscc_8924: i32_mulscc_Volatile port map(y_in => y_8544, A => operand_1_8671, B => operand_2_8677, Ni => Ni_8682, Zi => Zi_8687, Vi => Vi_8692, Ci => Ci_8697, y_out => i32_mulscc_y_8843, result => i32_mulscc_result_8843, No => Nmulscc_8843, Zo => Zmulscc_8843, Vo => Vmulscc_8843, Co => Cmulscc_8843); 
    volatile_operator_iu_umul32_8927: iu_umul32_Volatile port map(L => operand_1_8671, R => operand_2_8677, ret_val_x_x => uP_64_8853); 
    volatile_operator_i32_mul_calculate_sign_correction_8929: i32_mul_calculate_sign_correction_Volatile port map(signed_mul => signed_mul_div_8605, A => operand_1_8671, B => operand_2_8677, sign_correction => signed_correction_8862); 
    volatile_operator_exec_cti_instruction_8947: exec_cti_instruction_Volatile port map(exec_call => exec_call_8899, exec_rett => exec_rett_8905, exec_jmpl => exec_jmpl_8911, exec_ticc => exec_ticc_8917, br_cond => br_cond_8605, annul_flag => annul_flag_8605, pc => pc_8455, alu_result => i32_add_sub_result_8727, psr => psr_8516, wim => wim_8538, cti_trap_status => cti_trap_status_8951, cti_ticc_trap_type => cti_ticc_trap_type_8951, cti_trap_instr_trap => cti_trap_instr_trap_8951, cti_illegal_instr_trap => cti_illegal_instr_trap_8951, cti_privileged_instr_trap => cti_privileged_instr_trap_8951, cti_window_underflow_trap => cti_window_underflow_trap_8951, cti_mem_address_not_aligned_trap => cti_mem_address_not_aligned_trap_8951, cti_processor_error_mode => cti_processor_error_mode_8951, cti_br_taken => cti_br_taken_8951, cti_next_psr => cti_next_psr_8951, cti_annul_next => cti_annul_next_8951); 
    -- shared call operator group (9) : call_stmt_9223_call 
    i32_div_call_group_9: Block -- 
      signal data_in: std_logic_vector(97 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_9223_call_req_0;
      call_stmt_9223_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_9223_call_req_1;
      call_stmt_9223_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= issue_div_9211(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      i32_div_call_group_9_gI: SplitGuardInterface generic map(name => "i32_div_call_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= signed_mul_div_8605 & set_cc_8605 & y_8544 & operand_1_8671 & operand_2_8677;
      i32_div_result_9223 <= data_out(35 downto 4);
      Ndiv_9223 <= data_out(3 downto 3);
      Zdiv_9223 <= data_out(2 downto 2);
      Vdiv_9223 <= data_out(1 downto 1);
      Cdiv_9223 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 98,
        owidth => 98,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => i32_div_call_reqs(0),
          ackR => i32_div_call_acks(0),
          dataR => i32_div_call_data(97 downto 0),
          tagR => i32_div_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 36,
          owidth => 36,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => i32_div_return_acks(0), -- cross-over
          ackL => i32_div_return_reqs(0), -- cross-over
          dataL => i32_div_return_data(35 downto 0),
          tagL => i32_div_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 9
    -- 
  end Block; -- data_path
  -- 
end iu_exec_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity restore_window_trap_Volatile is -- 
  port ( -- 
    psr : in  std_logic_vector(31 downto 0);
    wim : in  std_logic_vector(31 downto 0);
    uflow_trap : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity restore_window_trap_Volatile;
architecture restore_window_trap_Volatile_arch of restore_window_trap_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(64-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal psr_buffer :  std_logic_vector(31 downto 0);
  signal wim_buffer :  std_logic_vector(31 downto 0);
  -- output port buffer signals
  signal uflow_trap_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  psr_buffer <= psr;
  wim_buffer <= wim;
  -- output handling  -------------------------------------------------------
  uflow_trap <= uflow_trap_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal ADD_u5_u5_8332_wire : std_logic_vector(4 downto 0);
    signal AND_u32_u32_8342_wire : std_logic_vector(31 downto 0);
    signal R_NWINDOWS_MOD_MASK_5_8333_wire_constant : std_logic_vector(4 downto 0);
    signal SHL_u32_u32_8341_wire : std_logic_vector(31 downto 0);
    signal curr_cwp_8328 : std_logic_vector(4 downto 0);
    signal konst_8331_wire_constant : std_logic_vector(4 downto 0);
    signal konst_8338_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8343_wire_constant : std_logic_vector(31 downto 0);
    signal new_cwp_8335 : std_logic_vector(4 downto 0);
    signal type_cast_8340_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_NWINDOWS_MOD_MASK_5_8333_wire_constant <= "00111";
    konst_8331_wire_constant <= "00001";
    konst_8338_wire_constant <= "00000000000000000000000000000001";
    konst_8343_wire_constant <= "00000000000000000000000000000000";
    -- flow-through slice operator slice_8327_inst
    curr_cwp_8328 <= psr_buffer(4 downto 0);
    -- interlock type_cast_8340_inst
    process(new_cwp_8335) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 4 downto 0) := new_cwp_8335(4 downto 0);
      type_cast_8340_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator ADD_u5_u5_8332_inst
    ADD_u5_u5_8332_wire <= std_logic_vector(unsigned(curr_cwp_8328) + unsigned(konst_8331_wire_constant));
    -- flow through binary operator AND_u32_u32_8342_inst
    AND_u32_u32_8342_wire <= (wim_buffer and SHL_u32_u32_8341_wire);
    -- flow through binary operator AND_u5_u5_8334_inst
    new_cwp_8335 <= (ADD_u5_u5_8332_wire and R_NWINDOWS_MOD_MASK_5_8333_wire_constant);
    -- flow through binary operator NEQ_u32_u1_8344_inst
    process(AND_u32_u32_8342_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(AND_u32_u32_8342_wire, konst_8343_wire_constant, tmp_var);
      uflow_trap_buffer <= tmp_var; --
    end process;
    -- flow through binary operator SHL_u32_u32_8341_inst
    process(konst_8338_wire_constant, type_cast_8340_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(konst_8338_wire_constant, type_cast_8340_wire, tmp_var);
      SHL_u32_u32_8341_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end restore_window_trap_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity save_window_trap_Volatile is -- 
  port ( -- 
    psr : in  std_logic_vector(31 downto 0);
    wim : in  std_logic_vector(31 downto 0);
    ovflow_trap : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity save_window_trap_Volatile;
architecture save_window_trap_Volatile_arch of save_window_trap_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(64-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal psr_buffer :  std_logic_vector(31 downto 0);
  signal wim_buffer :  std_logic_vector(31 downto 0);
  -- output port buffer signals
  signal ovflow_trap_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  psr_buffer <= psr;
  wim_buffer <= wim;
  -- output handling  -------------------------------------------------------
  ovflow_trap <= ovflow_trap_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u32_u32_8316_wire : std_logic_vector(31 downto 0);
    signal R_NWINDOWS_MOD_MASK_5_8307_wire_constant : std_logic_vector(4 downto 0);
    signal SHL_u32_u32_8315_wire : std_logic_vector(31 downto 0);
    signal SUB_u5_u5_8306_wire : std_logic_vector(4 downto 0);
    signal curr_cwp_8302 : std_logic_vector(4 downto 0);
    signal konst_8305_wire_constant : std_logic_vector(4 downto 0);
    signal konst_8312_wire_constant : std_logic_vector(31 downto 0);
    signal konst_8317_wire_constant : std_logic_vector(31 downto 0);
    signal new_cwp_8309 : std_logic_vector(4 downto 0);
    signal type_cast_8314_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_NWINDOWS_MOD_MASK_5_8307_wire_constant <= "00111";
    konst_8305_wire_constant <= "00001";
    konst_8312_wire_constant <= "00000000000000000000000000000001";
    konst_8317_wire_constant <= "00000000000000000000000000000000";
    -- flow-through slice operator slice_8301_inst
    curr_cwp_8302 <= psr_buffer(4 downto 0);
    -- interlock type_cast_8314_inst
    process(new_cwp_8309) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 4 downto 0) := new_cwp_8309(4 downto 0);
      type_cast_8314_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator AND_u32_u32_8316_inst
    AND_u32_u32_8316_wire <= (wim_buffer and SHL_u32_u32_8315_wire);
    -- flow through binary operator AND_u5_u5_8308_inst
    new_cwp_8309 <= (SUB_u5_u5_8306_wire and R_NWINDOWS_MOD_MASK_5_8307_wire_constant);
    -- flow through binary operator NEQ_u32_u1_8318_inst
    process(AND_u32_u32_8316_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(AND_u32_u32_8316_wire, konst_8317_wire_constant, tmp_var);
      ovflow_trap_buffer <= tmp_var; --
    end process;
    -- flow through binary operator SHL_u32_u32_8315_inst
    process(konst_8312_wire_constant, type_cast_8314_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(konst_8312_wire_constant, type_cast_8314_wire, tmp_var);
      SHL_u32_u32_8315_wire <= tmp_var; --
    end process;
    -- flow through binary operator SUB_u5_u5_8306_inst
    SUB_u5_u5_8306_wire <= std_logic_vector(unsigned(curr_cwp_8302) - unsigned(konst_8305_wire_constant));
    -- 
  end Block; -- data_path
  -- 
end save_window_trap_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity twos_complement_32_Volatile is -- 
  port ( -- 
    A : in  std_logic_vector(31 downto 0);
    B : out  std_logic_vector(31 downto 0)-- 
  );
  -- 
end entity twos_complement_32_Volatile;
architecture twos_complement_32_Volatile_arch of twos_complement_32_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(32-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal A_buffer :  std_logic_vector(31 downto 0);
  -- output port buffer signals
  signal B_buffer :  std_logic_vector(31 downto 0);
  -- volatile/operator module components. 
  component increment_32_Volatile is -- 
    port ( -- 
      A : in  std_logic_vector(31 downto 0);
      B : out  std_logic_vector(31 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  A_buffer <= A;
  -- output handling  -------------------------------------------------------
  B <= B_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal cA_7292 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    -- unary operator NOT_u32_u32_7291_inst
    process(A_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", A_buffer, tmp_var);
      cA_7292 <= tmp_var; -- 
    end process;
    volatile_operator_increment_32_6104: increment_32_Volatile port map(A => cA_7292, B => B_buffer); 
    -- 
  end Block; -- data_path
  -- 
end twos_complement_32_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity twos_complement_64_Volatile is -- 
  port ( -- 
    A : in  std_logic_vector(63 downto 0);
    B : out  std_logic_vector(63 downto 0)-- 
  );
  -- 
end entity twos_complement_64_Volatile;
architecture twos_complement_64_Volatile_arch of twos_complement_64_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(64-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal A_buffer :  std_logic_vector(63 downto 0);
  -- output port buffer signals
  signal B_buffer :  std_logic_vector(63 downto 0);
  -- volatile/operator module components. 
  component increment_64_Volatile is -- 
    port ( -- 
      A : in  std_logic_vector(63 downto 0);
      B : out  std_logic_vector(63 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  A_buffer <= A;
  -- output handling  -------------------------------------------------------
  B <= B_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal cA_7281 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    -- unary operator NOT_u64_u64_7280_inst
    process(A_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", A_buffer, tmp_var);
      cA_7281 <= tmp_var; -- 
    end process;
    volatile_operator_increment_64_6094: increment_64_Volatile port map(A => cA_7281, B => B_buffer); 
    -- 
  end Block; -- data_path
  -- 
end twos_complement_64_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity u32_sll_Volatile is -- 
  port ( -- 
    X : in  std_logic_vector(31 downto 0);
    S : in  std_logic_vector(5 downto 0);
    Y : out  std_logic_vector(31 downto 0)-- 
  );
  -- 
end entity u32_sll_Volatile;
architecture u32_sll_Volatile_arch of u32_sll_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(38-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal X_buffer :  std_logic_vector(31 downto 0);
  signal S_buffer :  std_logic_vector(5 downto 0);
  -- output port buffer signals
  signal Y_buffer :  std_logic_vector(31 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  X_buffer <= X;
  S_buffer <= S;
  -- output handling  -------------------------------------------------------
  Y <= Y_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u6_u1_1548_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u6_u1_1559_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u6_u1_1571_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u6_u1_1583_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u6_u1_1594_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u6_u1_1605_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u16_u32_1598_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u24_u32_1587_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u28_u32_1576_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u30_u32_1564_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u31_u32_1552_wire : std_logic_vector(31 downto 0);
    signal R_ZERO_16_1597_wire_constant : std_logic_vector(15 downto 0);
    signal R_ZERO_1_1551_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_2_1563_wire_constant : std_logic_vector(1 downto 0);
    signal R_ZERO_4_1575_wire_constant : std_logic_vector(3 downto 0);
    signal R_ZERO_8_1586_wire_constant : std_logic_vector(7 downto 0);
    signal X0_1555 : std_logic_vector(31 downto 0);
    signal X1_1567 : std_logic_vector(31 downto 0);
    signal X2_1579 : std_logic_vector(31 downto 0);
    signal X3_1590 : std_logic_vector(31 downto 0);
    signal X4_1601 : std_logic_vector(31 downto 0);
    signal konst_1547_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1558_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1570_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1582_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1593_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1604_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1606_wire_constant : std_logic_vector(31 downto 0);
    signal slice_1550_wire : std_logic_vector(30 downto 0);
    signal slice_1562_wire : std_logic_vector(29 downto 0);
    signal slice_1574_wire : std_logic_vector(27 downto 0);
    signal slice_1585_wire : std_logic_vector(23 downto 0);
    signal slice_1596_wire : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ZERO_16_1597_wire_constant <= "0000000000000000";
    R_ZERO_1_1551_wire_constant <= "0";
    R_ZERO_2_1563_wire_constant <= "00";
    R_ZERO_4_1575_wire_constant <= "0000";
    R_ZERO_8_1586_wire_constant <= "00000000";
    konst_1547_wire_constant <= "000000";
    konst_1558_wire_constant <= "000001";
    konst_1570_wire_constant <= "000010";
    konst_1582_wire_constant <= "000011";
    konst_1593_wire_constant <= "000100";
    konst_1604_wire_constant <= "000101";
    konst_1606_wire_constant <= "00000000000000000000000000000000";
    -- flow-through select operator MUX_1554_inst
    X0_1555 <= CONCAT_u31_u32_1552_wire when (BITSEL_u6_u1_1548_wire(0) /=  '0') else X_buffer;
    -- flow-through select operator MUX_1566_inst
    X1_1567 <= CONCAT_u30_u32_1564_wire when (BITSEL_u6_u1_1559_wire(0) /=  '0') else X0_1555;
    -- flow-through select operator MUX_1578_inst
    X2_1579 <= CONCAT_u28_u32_1576_wire when (BITSEL_u6_u1_1571_wire(0) /=  '0') else X1_1567;
    -- flow-through select operator MUX_1589_inst
    X3_1590 <= CONCAT_u24_u32_1587_wire when (BITSEL_u6_u1_1583_wire(0) /=  '0') else X2_1579;
    -- flow-through select operator MUX_1600_inst
    X4_1601 <= CONCAT_u16_u32_1598_wire when (BITSEL_u6_u1_1594_wire(0) /=  '0') else X3_1590;
    -- flow-through select operator MUX_1608_inst
    Y_buffer <= konst_1606_wire_constant when (BITSEL_u6_u1_1605_wire(0) /=  '0') else X4_1601;
    -- flow-through slice operator slice_1550_inst
    slice_1550_wire <= X_buffer(30 downto 0);
    -- flow-through slice operator slice_1562_inst
    slice_1562_wire <= X0_1555(29 downto 0);
    -- flow-through slice operator slice_1574_inst
    slice_1574_wire <= X1_1567(27 downto 0);
    -- flow-through slice operator slice_1585_inst
    slice_1585_wire <= X2_1579(23 downto 0);
    -- flow-through slice operator slice_1596_inst
    slice_1596_wire <= X3_1590(15 downto 0);
    -- flow through binary operator BITSEL_u6_u1_1548_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_1547_wire_constant, tmp_var);
      BITSEL_u6_u1_1548_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u6_u1_1559_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_1558_wire_constant, tmp_var);
      BITSEL_u6_u1_1559_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u6_u1_1571_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_1570_wire_constant, tmp_var);
      BITSEL_u6_u1_1571_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u6_u1_1583_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_1582_wire_constant, tmp_var);
      BITSEL_u6_u1_1583_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u6_u1_1594_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_1593_wire_constant, tmp_var);
      BITSEL_u6_u1_1594_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u6_u1_1605_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_1604_wire_constant, tmp_var);
      BITSEL_u6_u1_1605_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u16_u32_1598_inst
    process(slice_1596_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1596_wire, R_ZERO_16_1597_wire_constant, tmp_var);
      CONCAT_u16_u32_1598_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u24_u32_1587_inst
    process(slice_1585_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1585_wire, R_ZERO_8_1586_wire_constant, tmp_var);
      CONCAT_u24_u32_1587_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u28_u32_1576_inst
    process(slice_1574_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1574_wire, R_ZERO_4_1575_wire_constant, tmp_var);
      CONCAT_u28_u32_1576_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u30_u32_1564_inst
    process(slice_1562_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1562_wire, R_ZERO_2_1563_wire_constant, tmp_var);
      CONCAT_u30_u32_1564_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u31_u32_1552_inst
    process(slice_1550_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1550_wire, R_ZERO_1_1551_wire_constant, tmp_var);
      CONCAT_u31_u32_1552_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end u32_sll_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity u64_sll_Volatile is -- 
  port ( -- 
    X : in  std_logic_vector(63 downto 0);
    S : in  std_logic_vector(6 downto 0);
    Y : out  std_logic_vector(63 downto 0)-- 
  );
  -- 
end entity u64_sll_Volatile;
architecture u64_sll_Volatile_arch of u64_sll_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(71-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal X_buffer :  std_logic_vector(63 downto 0);
  signal S_buffer :  std_logic_vector(6 downto 0);
  -- output port buffer signals
  signal Y_buffer :  std_logic_vector(63 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  X_buffer <= X;
  S_buffer <= S;
  -- output handling  -------------------------------------------------------
  Y <= Y_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u7_u1_1467_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u7_u1_1478_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u7_u1_1489_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u7_u1_1501_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u7_u1_1513_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u7_u1_1524_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u7_u1_1535_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u32_u64_1528_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u48_u64_1517_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u56_u64_1506_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u60_u64_1494_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u62_u64_1482_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u63_u64_1471_wire : std_logic_vector(63 downto 0);
    signal R_ZERO_16_1516_wire_constant : std_logic_vector(15 downto 0);
    signal R_ZERO_1_1470_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_2_1481_wire_constant : std_logic_vector(1 downto 0);
    signal R_ZERO_32_1527_wire_constant : std_logic_vector(31 downto 0);
    signal R_ZERO_4_1493_wire_constant : std_logic_vector(3 downto 0);
    signal R_ZERO_8_1505_wire_constant : std_logic_vector(7 downto 0);
    signal X0_1474 : std_logic_vector(63 downto 0);
    signal X1_1485 : std_logic_vector(63 downto 0);
    signal X2_1497 : std_logic_vector(63 downto 0);
    signal X3_1509 : std_logic_vector(63 downto 0);
    signal X4_1520 : std_logic_vector(63 downto 0);
    signal X5_1531 : std_logic_vector(63 downto 0);
    signal konst_1466_wire_constant : std_logic_vector(6 downto 0);
    signal konst_1477_wire_constant : std_logic_vector(6 downto 0);
    signal konst_1488_wire_constant : std_logic_vector(6 downto 0);
    signal konst_1500_wire_constant : std_logic_vector(6 downto 0);
    signal konst_1512_wire_constant : std_logic_vector(6 downto 0);
    signal konst_1523_wire_constant : std_logic_vector(6 downto 0);
    signal konst_1534_wire_constant : std_logic_vector(6 downto 0);
    signal konst_1536_wire_constant : std_logic_vector(63 downto 0);
    signal slice_1469_wire : std_logic_vector(62 downto 0);
    signal slice_1480_wire : std_logic_vector(61 downto 0);
    signal slice_1492_wire : std_logic_vector(59 downto 0);
    signal slice_1504_wire : std_logic_vector(55 downto 0);
    signal slice_1515_wire : std_logic_vector(47 downto 0);
    signal slice_1526_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_ZERO_16_1516_wire_constant <= "0000000000000000";
    R_ZERO_1_1470_wire_constant <= "0";
    R_ZERO_2_1481_wire_constant <= "00";
    R_ZERO_32_1527_wire_constant <= "00000000000000000000000000000000";
    R_ZERO_4_1493_wire_constant <= "0000";
    R_ZERO_8_1505_wire_constant <= "00000000";
    konst_1466_wire_constant <= "0000000";
    konst_1477_wire_constant <= "0000001";
    konst_1488_wire_constant <= "0000010";
    konst_1500_wire_constant <= "0000011";
    konst_1512_wire_constant <= "0000100";
    konst_1523_wire_constant <= "0000101";
    konst_1534_wire_constant <= "0000110";
    konst_1536_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- flow-through select operator MUX_1473_inst
    X0_1474 <= CONCAT_u63_u64_1471_wire when (BITSEL_u7_u1_1467_wire(0) /=  '0') else X_buffer;
    -- flow-through select operator MUX_1484_inst
    X1_1485 <= CONCAT_u62_u64_1482_wire when (BITSEL_u7_u1_1478_wire(0) /=  '0') else X0_1474;
    -- flow-through select operator MUX_1496_inst
    X2_1497 <= CONCAT_u60_u64_1494_wire when (BITSEL_u7_u1_1489_wire(0) /=  '0') else X1_1485;
    -- flow-through select operator MUX_1508_inst
    X3_1509 <= CONCAT_u56_u64_1506_wire when (BITSEL_u7_u1_1501_wire(0) /=  '0') else X2_1497;
    -- flow-through select operator MUX_1519_inst
    X4_1520 <= CONCAT_u48_u64_1517_wire when (BITSEL_u7_u1_1513_wire(0) /=  '0') else X3_1509;
    -- flow-through select operator MUX_1530_inst
    X5_1531 <= CONCAT_u32_u64_1528_wire when (BITSEL_u7_u1_1524_wire(0) /=  '0') else X4_1520;
    -- flow-through select operator MUX_1538_inst
    Y_buffer <= konst_1536_wire_constant when (BITSEL_u7_u1_1535_wire(0) /=  '0') else X5_1531;
    -- flow-through slice operator slice_1469_inst
    slice_1469_wire <= X_buffer(62 downto 0);
    -- flow-through slice operator slice_1480_inst
    slice_1480_wire <= X0_1474(61 downto 0);
    -- flow-through slice operator slice_1492_inst
    slice_1492_wire <= X1_1485(59 downto 0);
    -- flow-through slice operator slice_1504_inst
    slice_1504_wire <= X2_1497(55 downto 0);
    -- flow-through slice operator slice_1515_inst
    slice_1515_wire <= X3_1509(47 downto 0);
    -- flow-through slice operator slice_1526_inst
    slice_1526_wire <= X4_1520(31 downto 0);
    -- flow through binary operator BITSEL_u7_u1_1467_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_1466_wire_constant, tmp_var);
      BITSEL_u7_u1_1467_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u7_u1_1478_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_1477_wire_constant, tmp_var);
      BITSEL_u7_u1_1478_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u7_u1_1489_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_1488_wire_constant, tmp_var);
      BITSEL_u7_u1_1489_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u7_u1_1501_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_1500_wire_constant, tmp_var);
      BITSEL_u7_u1_1501_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u7_u1_1513_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_1512_wire_constant, tmp_var);
      BITSEL_u7_u1_1513_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u7_u1_1524_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_1523_wire_constant, tmp_var);
      BITSEL_u7_u1_1524_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u7_u1_1535_inst
    process(S_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(S_buffer, konst_1534_wire_constant, tmp_var);
      BITSEL_u7_u1_1535_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u32_u64_1528_inst
    process(slice_1526_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1526_wire, R_ZERO_32_1527_wire_constant, tmp_var);
      CONCAT_u32_u64_1528_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u48_u64_1517_inst
    process(slice_1515_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1515_wire, R_ZERO_16_1516_wire_constant, tmp_var);
      CONCAT_u48_u64_1517_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u56_u64_1506_inst
    process(slice_1504_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1504_wire, R_ZERO_8_1505_wire_constant, tmp_var);
      CONCAT_u56_u64_1506_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u60_u64_1494_inst
    process(slice_1492_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1492_wire, R_ZERO_4_1493_wire_constant, tmp_var);
      CONCAT_u60_u64_1494_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u62_u64_1482_inst
    process(slice_1480_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1480_wire, R_ZERO_2_1481_wire_constant, tmp_var);
      CONCAT_u62_u64_1482_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u63_u64_1471_inst
    process(slice_1469_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1469_wire, R_ZERO_1_1470_wire_constant, tmp_var);
      CONCAT_u63_u64_1471_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end u64_sll_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity u64_true_divide_revised is -- 
  generic (tag_length : integer); 
  port ( -- 
    udividend : in  std_logic_vector(63 downto 0);
    udivisor : in  std_logic_vector(31 downto 0);
    quotient : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity u64_true_divide_revised;
architecture u64_true_divide_revised_arch of u64_true_divide_revised is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 96)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal udividend_buffer :  std_logic_vector(63 downto 0);
  signal udividend_update_enable: Boolean;
  signal udivisor_buffer :  std_logic_vector(31 downto 0);
  signal udivisor_update_enable: Boolean;
  -- output port buffer signals
  signal quotient_buffer :  std_logic_vector(63 downto 0);
  signal quotient_update_enable: Boolean;
  signal u64_true_divide_revised_CP_355_start: Boolean;
  signal u64_true_divide_revised_CP_355_symbol: Boolean;
  -- volatile/operator module components. 
  component alignDivisorToDividendRevised_Operator is -- 
    port ( -- 
      sample_req: in boolean;
      sample_ack: out boolean;
      update_req: in boolean;
      update_ack: out boolean;
      DIVIDEND : in  std_logic_vector(63 downto 0);
      udivisor : in  std_logic_vector(31 downto 0);
      SHIFTED_DIVIDEND : out  std_logic_vector(63 downto 0);
      SHIFTED_DIVISOR : out  std_logic_vector(31 downto 0);
      INITIAL_QMASK : out  std_logic_vector(63 downto 0);
      clk, reset: in std_logic
      -- 
    );
    -- 
  end component;
  component u64_true_divide_revised_core_Volatile is -- 
    port ( -- 
      QMASK : in  std_logic_vector(63 downto 0);
      QUOTIENT : in  std_logic_vector(63 downto 0);
      DIVIDEND : in  std_logic_vector(64 downto 0);
      SHIFTED_DIVISOR_34 : in  std_logic_vector(33 downto 0);
      SHIFTED_DIVISOR_34_2X : in  std_logic_vector(33 downto 0);
      SHIFTED_DIVISOR_34_3X : in  std_logic_vector(33 downto 0);
      COUNT : in  std_logic_vector(7 downto 0);
      NQMASK : out  std_logic_vector(63 downto 0);
      NQUOTIENT : out  std_logic_vector(63 downto 0);
      NDIVIDEND : out  std_logic_vector(64 downto 0);
      NCOUNT : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal phi_stmt_7510_req_1 : boolean;
  signal do_while_stmt_7508_branch_ack_0 : boolean;
  signal phi_stmt_7510_req_0 : boolean;
  signal do_while_stmt_7508_branch_req_0 : boolean;
  signal call_stmt_7489_call_ack_0 : boolean;
  signal call_stmt_7489_call_req_0 : boolean;
  signal INITIAL_QMASK_7489_7512_buf_ack_1 : boolean;
  signal NNQMASK_7567_7513_buf_req_0 : boolean;
  signal NNQMASK_7567_7513_buf_ack_0 : boolean;
  signal SHIFTED_DIVISOR_34_2X_7501_7539_buf_ack_0 : boolean;
  signal call_stmt_7489_call_req_1 : boolean;
  signal INITIAL_QMASK_7489_7512_buf_req_0 : boolean;
  signal INITIAL_QMASK_7489_7512_buf_req_1 : boolean;
  signal INITIAL_QMASK_7489_7512_buf_ack_0 : boolean;
  signal call_stmt_7489_call_ack_1 : boolean;
  signal phi_stmt_7510_ack_0 : boolean;
  signal NNQMASK_7567_7513_buf_ack_1 : boolean;
  signal NNQMASK_7567_7513_buf_req_1 : boolean;
  signal SHIFTED_DIVISOR_34_2X_7501_7539_buf_req_1 : boolean;
  signal phi_stmt_7514_req_1 : boolean;
  signal phi_stmt_7514_req_0 : boolean;
  signal phi_stmt_7514_ack_0 : boolean;
  signal NNQUOTIENT_7567_7517_buf_req_0 : boolean;
  signal NNQUOTIENT_7567_7517_buf_ack_0 : boolean;
  signal NNQUOTIENT_7567_7517_buf_req_1 : boolean;
  signal NNQUOTIENT_7567_7517_buf_ack_1 : boolean;
  signal phi_stmt_7518_req_0 : boolean;
  signal phi_stmt_7518_req_1 : boolean;
  signal phi_stmt_7518_ack_0 : boolean;
  signal NNDIVIDEND_7567_7520_buf_req_0 : boolean;
  signal NNDIVIDEND_7567_7520_buf_ack_0 : boolean;
  signal NNDIVIDEND_7567_7520_buf_req_1 : boolean;
  signal NNDIVIDEND_7567_7520_buf_ack_1 : boolean;
  signal CONCAT_u1_u65_7523_inst_req_0 : boolean;
  signal CONCAT_u1_u65_7523_inst_ack_0 : boolean;
  signal CONCAT_u1_u65_7523_inst_req_1 : boolean;
  signal CONCAT_u1_u65_7523_inst_ack_1 : boolean;
  signal phi_stmt_7524_req_1 : boolean;
  signal phi_stmt_7524_req_0 : boolean;
  signal phi_stmt_7524_ack_0 : boolean;
  signal SHIFTED_DIVISOR_34_2X_7501_7539_buf_ack_1 : boolean;
  signal NNCOUNT_7567_7527_buf_req_0 : boolean;
  signal NNCOUNT_7567_7527_buf_ack_0 : boolean;
  signal SHIFTED_DIVISOR_34_2X_7501_7539_buf_req_0 : boolean;
  signal NNCOUNT_7567_7527_buf_req_1 : boolean;
  signal NNCOUNT_7567_7527_buf_ack_1 : boolean;
  signal phi_stmt_7528_req_1 : boolean;
  signal phi_stmt_7528_req_0 : boolean;
  signal phi_stmt_7528_ack_0 : boolean;
  signal SHIFTED_DIVISOR_34_7496_7530_buf_req_0 : boolean;
  signal SHIFTED_DIVISOR_34_7496_7530_buf_ack_0 : boolean;
  signal do_while_stmt_7508_branch_ack_1 : boolean;
  signal SHIFTED_DIVISOR_34_7496_7530_buf_req_1 : boolean;
  signal SHIFTED_DIVISOR_34_7496_7530_buf_ack_1 : boolean;
  signal SHIFTED_DIVISOR_34_7496_7531_buf_req_0 : boolean;
  signal SHIFTED_DIVISOR_34_7496_7531_buf_ack_0 : boolean;
  signal SHIFTED_DIVISOR_34_7496_7531_buf_req_1 : boolean;
  signal SHIFTED_DIVISOR_34_7496_7531_buf_ack_1 : boolean;
  signal phi_stmt_7532_req_1 : boolean;
  signal phi_stmt_7532_req_0 : boolean;
  signal phi_stmt_7532_ack_0 : boolean;
  signal SHIFTED_DIVISOR_34_3X_7506_7534_buf_req_0 : boolean;
  signal SHIFTED_DIVISOR_34_3X_7506_7534_buf_ack_0 : boolean;
  signal SHIFTED_DIVISOR_34_3X_7506_7534_buf_req_1 : boolean;
  signal SHIFTED_DIVISOR_34_3X_7506_7534_buf_ack_1 : boolean;
  signal SHIFTED_DIVISOR_34_3X_7506_7535_buf_req_0 : boolean;
  signal SHIFTED_DIVISOR_34_3X_7506_7535_buf_ack_0 : boolean;
  signal SHIFTED_DIVISOR_34_3X_7506_7535_buf_req_1 : boolean;
  signal SHIFTED_DIVISOR_34_3X_7506_7535_buf_ack_1 : boolean;
  signal phi_stmt_7536_req_1 : boolean;
  signal phi_stmt_7536_req_0 : boolean;
  signal phi_stmt_7536_ack_0 : boolean;
  signal SHIFTED_DIVISOR_34_2X_7501_7538_buf_req_0 : boolean;
  signal SHIFTED_DIVISOR_34_2X_7501_7538_buf_ack_0 : boolean;
  signal SHIFTED_DIVISOR_34_2X_7501_7538_buf_req_1 : boolean;
  signal SHIFTED_DIVISOR_34_2X_7501_7538_buf_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "u64_true_divide_revised_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 96) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= udividend;
  udividend_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(95 downto 64) <= udivisor;
  udivisor_buffer <= in_buffer_data_out(95 downto 64);
  in_buffer_data_in(tag_length + 95 downto 96) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 95 downto 96);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  u64_true_divide_revised_CP_355_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "u64_true_divide_revised_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= quotient_buffer;
  quotient <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= u64_true_divide_revised_CP_355_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= u64_true_divide_revised_CP_355_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= u64_true_divide_revised_CP_355_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  u64_true_divide_revised_CP_355: Block -- control-path 
    signal u64_true_divide_revised_CP_355_elements: BooleanArray(154 downto 0);
    -- 
  begin -- 
    u64_true_divide_revised_CP_355_elements(0) <= u64_true_divide_revised_CP_355_start;
    u64_true_divide_revised_CP_355_symbol <= u64_true_divide_revised_CP_355_elements(3);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_7489_to_assign_stmt_7506/call_stmt_7489_Sample/$entry
      -- CP-element group 0: 	 call_stmt_7489_to_assign_stmt_7506/call_stmt_7489_Update/$entry
      -- CP-element group 0: 	 call_stmt_7489_to_assign_stmt_7506/call_stmt_7489_Sample/crr
      -- CP-element group 0: 	 call_stmt_7489_to_assign_stmt_7506/call_stmt_7489_Update/ccr
      -- CP-element group 0: 	 call_stmt_7489_to_assign_stmt_7506/call_stmt_7489_update_start_
      -- CP-element group 0: 	 call_stmt_7489_to_assign_stmt_7506/call_stmt_7489_sample_start_
      -- CP-element group 0: 	 call_stmt_7489_to_assign_stmt_7506/$entry
      -- CP-element group 0: 	 $entry
      -- 
    crr_368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(0), ack => call_stmt_7489_call_req_0); -- 
    ccr_373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(0), ack => call_stmt_7489_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_7489_to_assign_stmt_7506/call_stmt_7489_Sample/$exit
      -- CP-element group 1: 	 call_stmt_7489_to_assign_stmt_7506/call_stmt_7489_Sample/cra
      -- CP-element group 1: 	 call_stmt_7489_to_assign_stmt_7506/call_stmt_7489_sample_completed_
      -- 
    cra_369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_7489_call_ack_0, ack => u64_true_divide_revised_CP_355_elements(1)); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (7) 
      -- CP-element group 2: 	 call_stmt_7489_to_assign_stmt_7506/call_stmt_7489_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_7507/branch_block_stmt_7507__entry__
      -- CP-element group 2: 	 call_stmt_7489_to_assign_stmt_7506/call_stmt_7489_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_7507/do_while_stmt_7508__entry__
      -- CP-element group 2: 	 branch_block_stmt_7507/$entry
      -- CP-element group 2: 	 call_stmt_7489_to_assign_stmt_7506/call_stmt_7489_Update/cca
      -- CP-element group 2: 	 call_stmt_7489_to_assign_stmt_7506/$exit
      -- 
    cca_374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_7489_call_ack_1, ack => u64_true_divide_revised_CP_355_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	154 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_7507/do_while_stmt_7508__exit__
      -- CP-element group 3: 	 branch_block_stmt_7507/branch_block_stmt_7507__exit__
      -- CP-element group 3: 	 branch_block_stmt_7507/$exit
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 assign_stmt_7578/$exit
      -- CP-element group 3: 	 assign_stmt_7578/$entry
      -- 
    u64_true_divide_revised_CP_355_elements(3) <= u64_true_divide_revised_CP_355_elements(154);
    -- CP-element group 4:  transition  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_7507/do_while_stmt_7508/$entry
      -- CP-element group 4: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508__entry__
      -- 
    u64_true_divide_revised_CP_355_elements(4) <= u64_true_divide_revised_CP_355_elements(2);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	154 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508__exit__
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_7507/do_while_stmt_7508/loop_back
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	152 
    -- CP-element group 7: 	153 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_7507/do_while_stmt_7508/loop_exit/$entry
      -- CP-element group 7: 	 branch_block_stmt_7507/do_while_stmt_7508/condition_done
      -- CP-element group 7: 	 branch_block_stmt_7507/do_while_stmt_7508/loop_taken/$entry
      -- 
    u64_true_divide_revised_CP_355_elements(7) <= u64_true_divide_revised_CP_355_elements(12);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	14 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_7507/do_while_stmt_7508/loop_body_done
      -- 
    u64_true_divide_revised_CP_355_elements(8) <= u64_true_divide_revised_CP_355_elements(14);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	22 
    -- CP-element group 9: 	41 
    -- CP-element group 9: 	60 
    -- CP-element group 9: 	81 
    -- CP-element group 9: 	100 
    -- CP-element group 9: 	119 
    -- CP-element group 9: 	138 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/back_edge_to_loop_body
      -- 
    u64_true_divide_revised_CP_355_elements(9) <= u64_true_divide_revised_CP_355_elements(6);
    -- CP-element group 10:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	24 
    -- CP-element group 10: 	43 
    -- CP-element group 10: 	62 
    -- CP-element group 10: 	83 
    -- CP-element group 10: 	102 
    -- CP-element group 10: 	121 
    -- CP-element group 10: 	140 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/first_time_through_loop_body
      -- 
    u64_true_divide_revised_CP_355_elements(10) <= u64_true_divide_revised_CP_355_elements(4);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	19 
    -- CP-element group 11: 	35 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	54 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	75 
    -- CP-element group 11: 	76 
    -- CP-element group 11: 	94 
    -- CP-element group 11: 	95 
    -- CP-element group 11: 	113 
    -- CP-element group 11: 	114 
    -- CP-element group 11: 	132 
    -- CP-element group 11: 	133 
    -- CP-element group 11: 	151 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/$entry
      -- CP-element group 11: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/loop_body_start
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	21 
    -- CP-element group 12: 	40 
    -- CP-element group 12: 	59 
    -- CP-element group 12: 	80 
    -- CP-element group 12: 	99 
    -- CP-element group 12: 	118 
    -- CP-element group 12: 	137 
    -- CP-element group 12: 	151 
    -- CP-element group 12: 	15 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/condition_evaluated
      -- 
    condition_evaluated_396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(12), ack => do_while_stmt_7508_branch_req_0); -- 
    u64_true_divide_revised_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(17) & u64_true_divide_revised_CP_355_elements(21) & u64_true_divide_revised_CP_355_elements(40) & u64_true_divide_revised_CP_355_elements(59) & u64_true_divide_revised_CP_355_elements(80) & u64_true_divide_revised_CP_355_elements(99) & u64_true_divide_revised_CP_355_elements(118) & u64_true_divide_revised_CP_355_elements(137) & u64_true_divide_revised_CP_355_elements(151) & u64_true_divide_revised_CP_355_elements(15);
      gj_u64_true_divide_revised_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	18 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	54 
    -- CP-element group 13: 	75 
    -- CP-element group 13: 	94 
    -- CP-element group 13: 	113 
    -- CP-element group 13: 	132 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	17 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	37 
    -- CP-element group 13: 	56 
    -- CP-element group 13: 	77 
    -- CP-element group 13: 	96 
    -- CP-element group 13: 	115 
    -- CP-element group 13: 	134 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/aggregated_phi_sample_req
      -- CP-element group 13: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_sample_start__ps
      -- 
    u64_true_divide_revised_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(18) & u64_true_divide_revised_CP_355_elements(35) & u64_true_divide_revised_CP_355_elements(54) & u64_true_divide_revised_CP_355_elements(75) & u64_true_divide_revised_CP_355_elements(94) & u64_true_divide_revised_CP_355_elements(113) & u64_true_divide_revised_CP_355_elements(132) & u64_true_divide_revised_CP_355_elements(17);
      gj_u64_true_divide_revised_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	38 
    -- CP-element group 14: 	57 
    -- CP-element group 14: 	78 
    -- CP-element group 14: 	97 
    -- CP-element group 14: 	116 
    -- CP-element group 14: 	135 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	8 
    -- CP-element group 14: 	15 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	35 
    -- CP-element group 14: 	54 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	94 
    -- CP-element group 14: 	113 
    -- CP-element group 14: 	132 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/$exit
      -- CP-element group 14: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_sample_completed_
      -- 
    u64_true_divide_revised_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(20) & u64_true_divide_revised_CP_355_elements(38) & u64_true_divide_revised_CP_355_elements(57) & u64_true_divide_revised_CP_355_elements(78) & u64_true_divide_revised_CP_355_elements(97) & u64_true_divide_revised_CP_355_elements(116) & u64_true_divide_revised_CP_355_elements(135);
      gj_u64_true_divide_revised_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	12 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(15) is a control-delay.
    cp_element_15_delay: control_delay_element  generic map(name => " 15_delay", delay_value => 1)  port map(req => u64_true_divide_revised_CP_355_elements(14), ack => u64_true_divide_revised_CP_355_elements(15), clk => clk, reset =>reset);
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: 	36 
    -- CP-element group 16: 	55 
    -- CP-element group 16: 	76 
    -- CP-element group 16: 	95 
    -- CP-element group 16: 	114 
    -- CP-element group 16: 	133 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	39 
    -- CP-element group 16: 	58 
    -- CP-element group 16: 	79 
    -- CP-element group 16: 	98 
    -- CP-element group 16: 	117 
    -- CP-element group 16: 	136 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/aggregated_phi_update_req
      -- CP-element group 16: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_update_start__ps
      -- 
    u64_true_divide_revised_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(19) & u64_true_divide_revised_CP_355_elements(36) & u64_true_divide_revised_CP_355_elements(55) & u64_true_divide_revised_CP_355_elements(76) & u64_true_divide_revised_CP_355_elements(95) & u64_true_divide_revised_CP_355_elements(114) & u64_true_divide_revised_CP_355_elements(133);
      gj_u64_true_divide_revised_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	21 
    -- CP-element group 17: 	40 
    -- CP-element group 17: 	59 
    -- CP-element group 17: 	80 
    -- CP-element group 17: 	99 
    -- CP-element group 17: 	118 
    -- CP-element group 17: 	137 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/aggregated_phi_update_ack
      -- 
    u64_true_divide_revised_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(21) & u64_true_divide_revised_CP_355_elements(40) & u64_true_divide_revised_CP_355_elements(59) & u64_true_divide_revised_CP_355_elements(80) & u64_true_divide_revised_CP_355_elements(99) & u64_true_divide_revised_CP_355_elements(118) & u64_true_divide_revised_CP_355_elements(137);
      gj_u64_true_divide_revised_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	13 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_sample_start_
      -- 
    u64_true_divide_revised_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(14);
      gj_u64_true_divide_revised_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	11 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_update_start_
      -- 
    u64_true_divide_revised_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(21);
      gj_u64_true_divide_revised_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_sample_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: 	12 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_update_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	9 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_loopback_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(22) <= u64_true_divide_revised_CP_355_elements(9);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_loopback_sample_req
      -- CP-element group 23: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_loopback_sample_req_ps
      -- 
    phi_stmt_7510_loopback_sample_req_412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7510_loopback_sample_req_412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(23), ack => phi_stmt_7510_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	10 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_entry_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(24) <= u64_true_divide_revised_CP_355_elements(10);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_entry_sample_req_ps
      -- CP-element group 25: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_entry_sample_req
      -- 
    phi_stmt_7510_entry_sample_req_415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7510_entry_sample_req_415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(25), ack => phi_stmt_7510_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_phi_mux_ack_ps
      -- CP-element group 26: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7510_phi_mux_ack
      -- 
    phi_stmt_7510_phi_mux_ack_418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_7510_ack_0, ack => u64_true_divide_revised_CP_355_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_Sample/req
      -- CP-element group 27: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_sample_start__ps
      -- 
    req_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(27), ack => INITIAL_QMASK_7489_7512_buf_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_update_start__ps
      -- CP-element group 28: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_Update/req
      -- CP-element group 28: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_update_start_
      -- 
    req_436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(28), ack => INITIAL_QMASK_7489_7512_buf_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_Sample/ack
      -- CP-element group 29: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_sample_completed_
      -- 
    ack_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => INITIAL_QMASK_7489_7512_buf_ack_0, ack => u64_true_divide_revised_CP_355_elements(29)); -- 
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_Update/ack
      -- CP-element group 30: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_update_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_INITIAL_QMASK_7512_Update/$exit
      -- 
    ack_437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => INITIAL_QMASK_7489_7512_buf_ack_1, ack => u64_true_divide_revised_CP_355_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_Sample/req
      -- CP-element group 31: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_sample_start__ps
      -- 
    req_449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(31), ack => NNQMASK_7567_7513_buf_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_update_start_
      -- CP-element group 32: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_update_start__ps
      -- CP-element group 32: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_Update/req
      -- 
    req_454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(32), ack => NNQMASK_7567_7513_buf_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_sample_completed__ps
      -- 
    ack_450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NNQMASK_7567_7513_buf_ack_0, ack => u64_true_divide_revised_CP_355_elements(33)); -- 
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_Update/ack
      -- CP-element group 34: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQMASK_7513_update_completed__ps
      -- 
    ack_455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NNQMASK_7567_7513_buf_ack_1, ack => u64_true_divide_revised_CP_355_elements(34)); -- 
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	11 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	14 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_sample_start_
      -- 
    u64_true_divide_revised_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(14);
      gj_u64_true_divide_revised_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	40 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	16 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_update_start_
      -- 
    u64_true_divide_revised_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(40);
      gj_u64_true_divide_revised_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	13 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_sample_start__ps
      -- 
    u64_true_divide_revised_CP_355_elements(37) <= u64_true_divide_revised_CP_355_elements(13);
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	14 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_sample_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(38) is bound as output of CP function.
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	16 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_update_start__ps
      -- 
    u64_true_divide_revised_CP_355_elements(39) <= u64_true_divide_revised_CP_355_elements(16);
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	17 
    -- CP-element group 40: 	12 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	36 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_update_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	9 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_loopback_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(41) <= u64_true_divide_revised_CP_355_elements(9);
    -- CP-element group 42:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_loopback_sample_req
      -- CP-element group 42: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_loopback_sample_req_ps
      -- 
    phi_stmt_7514_loopback_sample_req_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7514_loopback_sample_req_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(42), ack => phi_stmt_7514_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	10 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_entry_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(43) <= u64_true_divide_revised_CP_355_elements(10);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_entry_sample_req
      -- CP-element group 44: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_entry_sample_req_ps
      -- 
    phi_stmt_7514_entry_sample_req_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7514_entry_sample_req_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(44), ack => phi_stmt_7514_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_phi_mux_ack
      -- CP-element group 45: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7514_phi_mux_ack_ps
      -- 
    phi_stmt_7514_phi_mux_ack_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_7514_ack_0, ack => u64_true_divide_revised_CP_355_elements(45)); -- 
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_64_7516_sample_start__ps
      -- CP-element group 46: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_64_7516_sample_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_64_7516_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_64_7516_sample_completed_
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_64_7516_update_start__ps
      -- CP-element group 47: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_64_7516_update_start_
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_64_7516_update_completed__ps
      -- 
    u64_true_divide_revised_CP_355_elements(48) <= u64_true_divide_revised_CP_355_elements(49);
    -- CP-element group 49:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	48 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_64_7516_update_completed_
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(49) is a control-delay.
    cp_element_49_delay: control_delay_element  generic map(name => " 49_delay", delay_value => 1)  port map(req => u64_true_divide_revised_CP_355_elements(47), ack => u64_true_divide_revised_CP_355_elements(49), clk => clk, reset =>reset);
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_sample_start__ps
      -- CP-element group 50: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_Sample/req
      -- 
    req_493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(50), ack => NNQUOTIENT_7567_7517_buf_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_update_start__ps
      -- CP-element group 51: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_update_start_
      -- CP-element group 51: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_Update/req
      -- 
    req_498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(51), ack => NNQUOTIENT_7567_7517_buf_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_sample_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_Sample/ack
      -- 
    ack_494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NNQUOTIENT_7567_7517_buf_ack_0, ack => u64_true_divide_revised_CP_355_elements(52)); -- 
    -- CP-element group 53:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_update_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNQUOTIENT_7517_Update/ack
      -- 
    ack_499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NNQUOTIENT_7567_7517_buf_ack_1, ack => u64_true_divide_revised_CP_355_elements(53)); -- 
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	11 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	14 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	13 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_sample_start_
      -- 
    u64_true_divide_revised_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(14);
      gj_u64_true_divide_revised_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	11 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	59 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	16 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_update_start_
      -- 
    u64_true_divide_revised_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(59);
      gj_u64_true_divide_revised_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	13 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_sample_start__ps
      -- 
    u64_true_divide_revised_CP_355_elements(56) <= u64_true_divide_revised_CP_355_elements(13);
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	14 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_sample_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(57) is bound as output of CP function.
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	16 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_update_start__ps
      -- 
    u64_true_divide_revised_CP_355_elements(58) <= u64_true_divide_revised_CP_355_elements(16);
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	17 
    -- CP-element group 59: 	12 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	55 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_update_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	9 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_loopback_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(60) <= u64_true_divide_revised_CP_355_elements(9);
    -- CP-element group 61:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_loopback_sample_req
      -- CP-element group 61: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_loopback_sample_req_ps
      -- 
    phi_stmt_7518_loopback_sample_req_510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7518_loopback_sample_req_510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(61), ack => phi_stmt_7518_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(61) is bound as output of CP function.
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	10 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_entry_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(62) <= u64_true_divide_revised_CP_355_elements(10);
    -- CP-element group 63:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_entry_sample_req
      -- CP-element group 63: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_entry_sample_req_ps
      -- 
    phi_stmt_7518_entry_sample_req_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7518_entry_sample_req_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(63), ack => phi_stmt_7518_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_phi_mux_ack
      -- CP-element group 64: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7518_phi_mux_ack_ps
      -- 
    phi_stmt_7518_phi_mux_ack_516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_7518_ack_0, ack => u64_true_divide_revised_CP_355_elements(64)); -- 
    -- CP-element group 65:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_sample_start__ps
      -- CP-element group 65: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_Sample/req
      -- 
    req_529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(65), ack => NNDIVIDEND_7567_7520_buf_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_update_start__ps
      -- CP-element group 66: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_update_start_
      -- CP-element group 66: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_Update/req
      -- 
    req_534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(66), ack => NNDIVIDEND_7567_7520_buf_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_sample_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_Sample/ack
      -- 
    ack_530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NNDIVIDEND_7567_7520_buf_ack_0, ack => u64_true_divide_revised_CP_355_elements(67)); -- 
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_update_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNDIVIDEND_7520_Update/ack
      -- 
    ack_535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NNDIVIDEND_7567_7520_buf_ack_1, ack => u64_true_divide_revised_CP_355_elements(68)); -- 
    -- CP-element group 69:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_sample_start__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_update_start__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_Sample/rr
      -- 
    rr_547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(71), ack => CONCAT_u1_u65_7523_inst_req_0); -- 
    u64_true_divide_revised_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(69) & u64_true_divide_revised_CP_355_elements(73);
      gj_u64_true_divide_revised_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	74 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_update_start_
      -- CP-element group 72: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_Update/cr
      -- 
    cr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(72), ack => CONCAT_u1_u65_7523_inst_req_1); -- 
    u64_true_divide_revised_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(70) & u64_true_divide_revised_CP_355_elements(74);
      gj_u64_true_divide_revised_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_sample_completed__ps
      -- CP-element group 73: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_Sample/ra
      -- 
    ra_548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u65_7523_inst_ack_0, ack => u64_true_divide_revised_CP_355_elements(73)); -- 
    -- CP-element group 74:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	72 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_update_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/CONCAT_u1_u65_7523_Update/ca
      -- 
    ca_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u65_7523_inst_ack_1, ack => u64_true_divide_revised_CP_355_elements(74)); -- 
    -- CP-element group 75:  join  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	11 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	13 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_sample_start_
      -- 
    u64_true_divide_revised_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(14);
      gj_u64_true_divide_revised_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	11 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	80 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	16 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_update_start_
      -- 
    u64_true_divide_revised_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(80);
      gj_u64_true_divide_revised_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	13 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_sample_start__ps
      -- 
    u64_true_divide_revised_CP_355_elements(77) <= u64_true_divide_revised_CP_355_elements(13);
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	14 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_sample_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(78) is bound as output of CP function.
    -- CP-element group 79:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	16 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_update_start__ps
      -- 
    u64_true_divide_revised_CP_355_elements(79) <= u64_true_divide_revised_CP_355_elements(16);
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	17 
    -- CP-element group 80: 	12 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	76 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_update_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(80) is bound as output of CP function.
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	9 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_loopback_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(81) <= u64_true_divide_revised_CP_355_elements(9);
    -- CP-element group 82:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_loopback_sample_req
      -- CP-element group 82: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_loopback_sample_req_ps
      -- 
    phi_stmt_7524_loopback_sample_req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7524_loopback_sample_req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(82), ack => phi_stmt_7524_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(82) is bound as output of CP function.
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	10 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_entry_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(83) <= u64_true_divide_revised_CP_355_elements(10);
    -- CP-element group 84:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_entry_sample_req
      -- CP-element group 84: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_entry_sample_req_ps
      -- 
    phi_stmt_7524_entry_sample_req_567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7524_entry_sample_req_567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(84), ack => phi_stmt_7524_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(84) is bound as output of CP function.
    -- CP-element group 85:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_phi_mux_ack
      -- CP-element group 85: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7524_phi_mux_ack_ps
      -- 
    phi_stmt_7524_phi_mux_ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_7524_ack_0, ack => u64_true_divide_revised_CP_355_elements(85)); -- 
    -- CP-element group 86:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_8_7526_sample_start__ps
      -- CP-element group 86: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_8_7526_sample_completed__ps
      -- CP-element group 86: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_8_7526_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_8_7526_sample_completed_
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_8_7526_update_start__ps
      -- CP-element group 87: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_8_7526_update_start_
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_8_7526_update_completed__ps
      -- 
    u64_true_divide_revised_CP_355_elements(88) <= u64_true_divide_revised_CP_355_elements(89);
    -- CP-element group 89:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	88 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_ZERO_8_7526_update_completed_
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => u64_true_divide_revised_CP_355_elements(87), ack => u64_true_divide_revised_CP_355_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_sample_start__ps
      -- CP-element group 90: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_Sample/req
      -- 
    req_591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(90), ack => NNCOUNT_7567_7527_buf_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_update_start__ps
      -- CP-element group 91: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_update_start_
      -- CP-element group 91: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_Update/req
      -- 
    req_596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(91), ack => NNCOUNT_7567_7527_buf_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(91) is bound as output of CP function.
    -- CP-element group 92:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (4) 
      -- CP-element group 92: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_sample_completed__ps
      -- CP-element group 92: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_Sample/ack
      -- 
    ack_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NNCOUNT_7567_7527_buf_ack_0, ack => u64_true_divide_revised_CP_355_elements(92)); -- 
    -- CP-element group 93:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_update_completed__ps
      -- CP-element group 93: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_NNCOUNT_7527_Update/ack
      -- 
    ack_597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NNCOUNT_7567_7527_buf_ack_1, ack => u64_true_divide_revised_CP_355_elements(93)); -- 
    -- CP-element group 94:  join  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	11 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	14 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	13 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_sample_start_
      -- 
    u64_true_divide_revised_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(14);
      gj_u64_true_divide_revised_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	11 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	99 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	16 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_update_start_
      -- 
    u64_true_divide_revised_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "u64_true_divide_revised_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(99);
      gj_u64_true_divide_revised_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	13 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_sample_start__ps
      -- 
    u64_true_divide_revised_CP_355_elements(96) <= u64_true_divide_revised_CP_355_elements(13);
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	14 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_sample_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(97) is bound as output of CP function.
    -- CP-element group 98:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	16 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_update_start__ps
      -- 
    u64_true_divide_revised_CP_355_elements(98) <= u64_true_divide_revised_CP_355_elements(16);
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	17 
    -- CP-element group 99: 	12 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	95 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_update_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(99) is bound as output of CP function.
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	9 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_loopback_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(100) <= u64_true_divide_revised_CP_355_elements(9);
    -- CP-element group 101:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_loopback_sample_req
      -- CP-element group 101: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_loopback_sample_req_ps
      -- 
    phi_stmt_7528_loopback_sample_req_608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7528_loopback_sample_req_608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(101), ack => phi_stmt_7528_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(101) is bound as output of CP function.
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	10 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_entry_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(102) <= u64_true_divide_revised_CP_355_elements(10);
    -- CP-element group 103:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_entry_sample_req
      -- CP-element group 103: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_entry_sample_req_ps
      -- 
    phi_stmt_7528_entry_sample_req_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7528_entry_sample_req_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(103), ack => phi_stmt_7528_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(103) is bound as output of CP function.
    -- CP-element group 104:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_phi_mux_ack
      -- CP-element group 104: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7528_phi_mux_ack_ps
      -- 
    phi_stmt_7528_phi_mux_ack_614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_7528_ack_0, ack => u64_true_divide_revised_CP_355_elements(104)); -- 
    -- CP-element group 105:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_sample_start__ps
      -- CP-element group 105: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_Sample/req
      -- 
    req_627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(105), ack => SHIFTED_DIVISOR_34_7496_7530_buf_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_update_start__ps
      -- CP-element group 106: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_update_start_
      -- CP-element group 106: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_Update/req
      -- 
    req_632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(106), ack => SHIFTED_DIVISOR_34_7496_7530_buf_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_sample_completed__ps
      -- CP-element group 107: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_Sample/ack
      -- 
    ack_628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHIFTED_DIVISOR_34_7496_7530_buf_ack_0, ack => u64_true_divide_revised_CP_355_elements(107)); -- 
    -- CP-element group 108:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_update_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7530_Update/ack
      -- 
    ack_633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHIFTED_DIVISOR_34_7496_7530_buf_ack_1, ack => u64_true_divide_revised_CP_355_elements(108)); -- 
    -- CP-element group 109:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_sample_start__ps
      -- CP-element group 109: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_Sample/req
      -- 
    req_645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(109), ack => SHIFTED_DIVISOR_34_7496_7531_buf_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (4) 
      -- CP-element group 110: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_update_start__ps
      -- CP-element group 110: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_update_start_
      -- CP-element group 110: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_Update/req
      -- 
    req_650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(110), ack => SHIFTED_DIVISOR_34_7496_7531_buf_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(110) is bound as output of CP function.
    -- CP-element group 111:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (4) 
      -- CP-element group 111: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_sample_completed__ps
      -- CP-element group 111: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_Sample/ack
      -- 
    ack_646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHIFTED_DIVISOR_34_7496_7531_buf_ack_0, ack => u64_true_divide_revised_CP_355_elements(111)); -- 
    -- CP-element group 112:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_update_completed__ps
      -- CP-element group 112: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_7531_Update/ack
      -- 
    ack_651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHIFTED_DIVISOR_34_7496_7531_buf_ack_1, ack => u64_true_divide_revised_CP_355_elements(112)); -- 
    -- CP-element group 113:  join  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	11 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	14 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	13 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_sample_start_
      -- 
    u64_true_divide_revised_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "u64_true_divide_revised_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(14);
      gj_u64_true_divide_revised_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	11 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	118 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	16 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_update_start_
      -- 
    u64_true_divide_revised_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "u64_true_divide_revised_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(118);
      gj_u64_true_divide_revised_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	13 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_sample_start__ps
      -- 
    u64_true_divide_revised_CP_355_elements(115) <= u64_true_divide_revised_CP_355_elements(13);
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	14 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_sample_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(116) is bound as output of CP function.
    -- CP-element group 117:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	16 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_update_start__ps
      -- 
    u64_true_divide_revised_CP_355_elements(117) <= u64_true_divide_revised_CP_355_elements(16);
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	17 
    -- CP-element group 118: 	12 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	114 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_update_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(118) is bound as output of CP function.
    -- CP-element group 119:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	9 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_loopback_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(119) <= u64_true_divide_revised_CP_355_elements(9);
    -- CP-element group 120:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_loopback_sample_req
      -- CP-element group 120: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_loopback_sample_req_ps
      -- 
    phi_stmt_7532_loopback_sample_req_662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7532_loopback_sample_req_662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(120), ack => phi_stmt_7532_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(120) is bound as output of CP function.
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	10 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_entry_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(121) <= u64_true_divide_revised_CP_355_elements(10);
    -- CP-element group 122:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_entry_sample_req
      -- CP-element group 122: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_entry_sample_req_ps
      -- 
    phi_stmt_7532_entry_sample_req_665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7532_entry_sample_req_665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(122), ack => phi_stmt_7532_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(122) is bound as output of CP function.
    -- CP-element group 123:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_phi_mux_ack
      -- CP-element group 123: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7532_phi_mux_ack_ps
      -- 
    phi_stmt_7532_phi_mux_ack_668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_7532_ack_0, ack => u64_true_divide_revised_CP_355_elements(123)); -- 
    -- CP-element group 124:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (4) 
      -- CP-element group 124: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_sample_start__ps
      -- CP-element group 124: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_Sample/req
      -- 
    req_681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(124), ack => SHIFTED_DIVISOR_34_3X_7506_7534_buf_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(124) is bound as output of CP function.
    -- CP-element group 125:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_update_start__ps
      -- CP-element group 125: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_update_start_
      -- CP-element group 125: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_Update/$entry
      -- CP-element group 125: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_Update/req
      -- 
    req_686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(125), ack => SHIFTED_DIVISOR_34_3X_7506_7534_buf_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_sample_completed__ps
      -- CP-element group 126: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_Sample/ack
      -- 
    ack_682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHIFTED_DIVISOR_34_3X_7506_7534_buf_ack_0, ack => u64_true_divide_revised_CP_355_elements(126)); -- 
    -- CP-element group 127:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_update_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7534_Update/ack
      -- 
    ack_687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHIFTED_DIVISOR_34_3X_7506_7534_buf_ack_1, ack => u64_true_divide_revised_CP_355_elements(127)); -- 
    -- CP-element group 128:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (4) 
      -- CP-element group 128: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_sample_start__ps
      -- CP-element group 128: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_Sample/req
      -- 
    req_699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(128), ack => SHIFTED_DIVISOR_34_3X_7506_7535_buf_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (4) 
      -- CP-element group 129: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_update_start__ps
      -- CP-element group 129: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_update_start_
      -- CP-element group 129: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_Update/req
      -- 
    req_704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(129), ack => SHIFTED_DIVISOR_34_3X_7506_7535_buf_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (4) 
      -- CP-element group 130: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_sample_completed__ps
      -- CP-element group 130: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_Sample/ack
      -- 
    ack_700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHIFTED_DIVISOR_34_3X_7506_7535_buf_ack_0, ack => u64_true_divide_revised_CP_355_elements(130)); -- 
    -- CP-element group 131:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (4) 
      -- CP-element group 131: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_update_completed__ps
      -- CP-element group 131: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_3X_7535_Update/ack
      -- 
    ack_705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHIFTED_DIVISOR_34_3X_7506_7535_buf_ack_1, ack => u64_true_divide_revised_CP_355_elements(131)); -- 
    -- CP-element group 132:  join  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	11 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	14 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	13 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_sample_start_
      -- 
    u64_true_divide_revised_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "u64_true_divide_revised_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(14);
      gj_u64_true_divide_revised_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	11 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	137 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	16 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_update_start_
      -- 
    u64_true_divide_revised_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "u64_true_divide_revised_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= u64_true_divide_revised_CP_355_elements(11) & u64_true_divide_revised_CP_355_elements(137);
      gj_u64_true_divide_revised_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	13 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_sample_start__ps
      -- 
    u64_true_divide_revised_CP_355_elements(134) <= u64_true_divide_revised_CP_355_elements(13);
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	14 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_sample_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(135) is bound as output of CP function.
    -- CP-element group 136:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	16 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_update_start__ps
      -- 
    u64_true_divide_revised_CP_355_elements(136) <= u64_true_divide_revised_CP_355_elements(16);
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	17 
    -- CP-element group 137: 	12 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	133 
    -- CP-element group 137:  members (2) 
      -- CP-element group 137: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_update_completed__ps
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(137) is bound as output of CP function.
    -- CP-element group 138:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	9 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_loopback_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(138) <= u64_true_divide_revised_CP_355_elements(9);
    -- CP-element group 139:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (2) 
      -- CP-element group 139: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_loopback_sample_req
      -- CP-element group 139: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_loopback_sample_req_ps
      -- 
    phi_stmt_7536_loopback_sample_req_716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7536_loopback_sample_req_716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(139), ack => phi_stmt_7536_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(139) is bound as output of CP function.
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	10 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_entry_trigger
      -- 
    u64_true_divide_revised_CP_355_elements(140) <= u64_true_divide_revised_CP_355_elements(10);
    -- CP-element group 141:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_entry_sample_req
      -- CP-element group 141: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_entry_sample_req_ps
      -- 
    phi_stmt_7536_entry_sample_req_719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_7536_entry_sample_req_719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(141), ack => phi_stmt_7536_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(141) is bound as output of CP function.
    -- CP-element group 142:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_phi_mux_ack
      -- CP-element group 142: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/phi_stmt_7536_phi_mux_ack_ps
      -- 
    phi_stmt_7536_phi_mux_ack_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_7536_ack_0, ack => u64_true_divide_revised_CP_355_elements(142)); -- 
    -- CP-element group 143:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (4) 
      -- CP-element group 143: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_sample_start__ps
      -- CP-element group 143: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_Sample/req
      -- 
    req_735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(143), ack => SHIFTED_DIVISOR_34_2X_7501_7538_buf_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(143) is bound as output of CP function.
    -- CP-element group 144:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_update_start__ps
      -- CP-element group 144: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_update_start_
      -- CP-element group 144: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_Update/req
      -- 
    req_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(144), ack => SHIFTED_DIVISOR_34_2X_7501_7538_buf_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (4) 
      -- CP-element group 145: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_sample_completed__ps
      -- CP-element group 145: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_Sample/ack
      -- 
    ack_736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHIFTED_DIVISOR_34_2X_7501_7538_buf_ack_0, ack => u64_true_divide_revised_CP_355_elements(145)); -- 
    -- CP-element group 146:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_update_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7538_Update/ack
      -- 
    ack_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHIFTED_DIVISOR_34_2X_7501_7538_buf_ack_1, ack => u64_true_divide_revised_CP_355_elements(146)); -- 
    -- CP-element group 147:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (4) 
      -- CP-element group 147: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_Sample/req
      -- CP-element group 147: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_sample_start__ps
      -- 
    req_753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(147), ack => SHIFTED_DIVISOR_34_2X_7501_7539_buf_req_0); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (4) 
      -- CP-element group 148: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_update_start_
      -- CP-element group 148: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_Update/req
      -- CP-element group 148: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_update_start__ps
      -- 
    req_758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => u64_true_divide_revised_CP_355_elements(148), ack => SHIFTED_DIVISOR_34_2X_7501_7539_buf_req_1); -- 
    -- Element group u64_true_divide_revised_CP_355_elements(148) is bound as output of CP function.
    -- CP-element group 149:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (4) 
      -- CP-element group 149: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_Sample/ack
      -- CP-element group 149: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_sample_completed__ps
      -- 
    ack_754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHIFTED_DIVISOR_34_2X_7501_7539_buf_ack_0, ack => u64_true_divide_revised_CP_355_elements(149)); -- 
    -- CP-element group 150:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_Update/ack
      -- CP-element group 150: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/R_SHIFTED_DIVISOR_34_2X_7539_update_completed__ps
      -- 
    ack_759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHIFTED_DIVISOR_34_2X_7501_7539_buf_ack_1, ack => u64_true_divide_revised_CP_355_elements(150)); -- 
    -- CP-element group 151:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	11 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	12 
    -- CP-element group 151:  members (1) 
      -- CP-element group 151: 	 branch_block_stmt_7507/do_while_stmt_7508/do_while_stmt_7508_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group u64_true_divide_revised_CP_355_elements(151) is a control-delay.
    cp_element_151_delay: control_delay_element  generic map(name => " 151_delay", delay_value => 1)  port map(req => u64_true_divide_revised_CP_355_elements(11), ack => u64_true_divide_revised_CP_355_elements(151), clk => clk, reset =>reset);
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	7 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (2) 
      -- CP-element group 152: 	 branch_block_stmt_7507/do_while_stmt_7508/loop_exit/ack
      -- CP-element group 152: 	 branch_block_stmt_7507/do_while_stmt_7508/loop_exit/$exit
      -- 
    ack_765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_7508_branch_ack_0, ack => u64_true_divide_revised_CP_355_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	7 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (2) 
      -- CP-element group 153: 	 branch_block_stmt_7507/do_while_stmt_7508/loop_taken/ack
      -- CP-element group 153: 	 branch_block_stmt_7507/do_while_stmt_7508/loop_taken/$exit
      -- 
    ack_769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_7508_branch_ack_1, ack => u64_true_divide_revised_CP_355_elements(153)); -- 
    -- CP-element group 154:  transition  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	5 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	3 
    -- CP-element group 154:  members (1) 
      -- CP-element group 154: 	 branch_block_stmt_7507/do_while_stmt_7508/$exit
      -- 
    u64_true_divide_revised_CP_355_elements(154) <= u64_true_divide_revised_CP_355_elements(5);
    u64_true_divide_revised_do_while_stmt_7508_terminator_770: loop_terminator -- 
      generic map (name => " u64_true_divide_revised_do_while_stmt_7508_terminator_770", max_iterations_in_flight =>7) 
      port map(loop_body_exit => u64_true_divide_revised_CP_355_elements(8),loop_continue => u64_true_divide_revised_CP_355_elements(153),loop_terminate => u64_true_divide_revised_CP_355_elements(152),loop_back => u64_true_divide_revised_CP_355_elements(6),loop_exit => u64_true_divide_revised_CP_355_elements(5),clk => clk, reset => reset); -- 
    phi_stmt_7510_phi_seq_456_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= u64_true_divide_revised_CP_355_elements(24);
      u64_true_divide_revised_CP_355_elements(27)<= src_sample_reqs(0);
      src_sample_acks(0)  <= u64_true_divide_revised_CP_355_elements(29);
      u64_true_divide_revised_CP_355_elements(28)<= src_update_reqs(0);
      src_update_acks(0)  <= u64_true_divide_revised_CP_355_elements(30);
      u64_true_divide_revised_CP_355_elements(25) <= phi_mux_reqs(0);
      triggers(1)  <= u64_true_divide_revised_CP_355_elements(22);
      u64_true_divide_revised_CP_355_elements(31)<= src_sample_reqs(1);
      src_sample_acks(1)  <= u64_true_divide_revised_CP_355_elements(33);
      u64_true_divide_revised_CP_355_elements(32)<= src_update_reqs(1);
      src_update_acks(1)  <= u64_true_divide_revised_CP_355_elements(34);
      u64_true_divide_revised_CP_355_elements(23) <= phi_mux_reqs(1);
      phi_stmt_7510_phi_seq_456 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_7510_phi_seq_456") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => u64_true_divide_revised_CP_355_elements(13), 
          phi_sample_ack => u64_true_divide_revised_CP_355_elements(20), 
          phi_update_req => u64_true_divide_revised_CP_355_elements(16), 
          phi_update_ack => u64_true_divide_revised_CP_355_elements(21), 
          phi_mux_ack => u64_true_divide_revised_CP_355_elements(26), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_7514_phi_seq_500_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= u64_true_divide_revised_CP_355_elements(43);
      u64_true_divide_revised_CP_355_elements(46)<= src_sample_reqs(0);
      src_sample_acks(0)  <= u64_true_divide_revised_CP_355_elements(46);
      u64_true_divide_revised_CP_355_elements(47)<= src_update_reqs(0);
      src_update_acks(0)  <= u64_true_divide_revised_CP_355_elements(48);
      u64_true_divide_revised_CP_355_elements(44) <= phi_mux_reqs(0);
      triggers(1)  <= u64_true_divide_revised_CP_355_elements(41);
      u64_true_divide_revised_CP_355_elements(50)<= src_sample_reqs(1);
      src_sample_acks(1)  <= u64_true_divide_revised_CP_355_elements(52);
      u64_true_divide_revised_CP_355_elements(51)<= src_update_reqs(1);
      src_update_acks(1)  <= u64_true_divide_revised_CP_355_elements(53);
      u64_true_divide_revised_CP_355_elements(42) <= phi_mux_reqs(1);
      phi_stmt_7514_phi_seq_500 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_7514_phi_seq_500") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => u64_true_divide_revised_CP_355_elements(37), 
          phi_sample_ack => u64_true_divide_revised_CP_355_elements(38), 
          phi_update_req => u64_true_divide_revised_CP_355_elements(39), 
          phi_update_ack => u64_true_divide_revised_CP_355_elements(40), 
          phi_mux_ack => u64_true_divide_revised_CP_355_elements(45), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_7518_phi_seq_554_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= u64_true_divide_revised_CP_355_elements(60);
      u64_true_divide_revised_CP_355_elements(65)<= src_sample_reqs(0);
      src_sample_acks(0)  <= u64_true_divide_revised_CP_355_elements(67);
      u64_true_divide_revised_CP_355_elements(66)<= src_update_reqs(0);
      src_update_acks(0)  <= u64_true_divide_revised_CP_355_elements(68);
      u64_true_divide_revised_CP_355_elements(61) <= phi_mux_reqs(0);
      triggers(1)  <= u64_true_divide_revised_CP_355_elements(62);
      u64_true_divide_revised_CP_355_elements(69)<= src_sample_reqs(1);
      src_sample_acks(1)  <= u64_true_divide_revised_CP_355_elements(73);
      u64_true_divide_revised_CP_355_elements(70)<= src_update_reqs(1);
      src_update_acks(1)  <= u64_true_divide_revised_CP_355_elements(74);
      u64_true_divide_revised_CP_355_elements(63) <= phi_mux_reqs(1);
      phi_stmt_7518_phi_seq_554 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_7518_phi_seq_554") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => u64_true_divide_revised_CP_355_elements(56), 
          phi_sample_ack => u64_true_divide_revised_CP_355_elements(57), 
          phi_update_req => u64_true_divide_revised_CP_355_elements(58), 
          phi_update_ack => u64_true_divide_revised_CP_355_elements(59), 
          phi_mux_ack => u64_true_divide_revised_CP_355_elements(64), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_7524_phi_seq_598_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= u64_true_divide_revised_CP_355_elements(83);
      u64_true_divide_revised_CP_355_elements(86)<= src_sample_reqs(0);
      src_sample_acks(0)  <= u64_true_divide_revised_CP_355_elements(86);
      u64_true_divide_revised_CP_355_elements(87)<= src_update_reqs(0);
      src_update_acks(0)  <= u64_true_divide_revised_CP_355_elements(88);
      u64_true_divide_revised_CP_355_elements(84) <= phi_mux_reqs(0);
      triggers(1)  <= u64_true_divide_revised_CP_355_elements(81);
      u64_true_divide_revised_CP_355_elements(90)<= src_sample_reqs(1);
      src_sample_acks(1)  <= u64_true_divide_revised_CP_355_elements(92);
      u64_true_divide_revised_CP_355_elements(91)<= src_update_reqs(1);
      src_update_acks(1)  <= u64_true_divide_revised_CP_355_elements(93);
      u64_true_divide_revised_CP_355_elements(82) <= phi_mux_reqs(1);
      phi_stmt_7524_phi_seq_598 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_7524_phi_seq_598") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => u64_true_divide_revised_CP_355_elements(77), 
          phi_sample_ack => u64_true_divide_revised_CP_355_elements(78), 
          phi_update_req => u64_true_divide_revised_CP_355_elements(79), 
          phi_update_ack => u64_true_divide_revised_CP_355_elements(80), 
          phi_mux_ack => u64_true_divide_revised_CP_355_elements(85), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_7528_phi_seq_652_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= u64_true_divide_revised_CP_355_elements(102);
      u64_true_divide_revised_CP_355_elements(105)<= src_sample_reqs(0);
      src_sample_acks(0)  <= u64_true_divide_revised_CP_355_elements(107);
      u64_true_divide_revised_CP_355_elements(106)<= src_update_reqs(0);
      src_update_acks(0)  <= u64_true_divide_revised_CP_355_elements(108);
      u64_true_divide_revised_CP_355_elements(103) <= phi_mux_reqs(0);
      triggers(1)  <= u64_true_divide_revised_CP_355_elements(100);
      u64_true_divide_revised_CP_355_elements(109)<= src_sample_reqs(1);
      src_sample_acks(1)  <= u64_true_divide_revised_CP_355_elements(111);
      u64_true_divide_revised_CP_355_elements(110)<= src_update_reqs(1);
      src_update_acks(1)  <= u64_true_divide_revised_CP_355_elements(112);
      u64_true_divide_revised_CP_355_elements(101) <= phi_mux_reqs(1);
      phi_stmt_7528_phi_seq_652 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_7528_phi_seq_652") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => u64_true_divide_revised_CP_355_elements(96), 
          phi_sample_ack => u64_true_divide_revised_CP_355_elements(97), 
          phi_update_req => u64_true_divide_revised_CP_355_elements(98), 
          phi_update_ack => u64_true_divide_revised_CP_355_elements(99), 
          phi_mux_ack => u64_true_divide_revised_CP_355_elements(104), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_7532_phi_seq_706_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= u64_true_divide_revised_CP_355_elements(121);
      u64_true_divide_revised_CP_355_elements(124)<= src_sample_reqs(0);
      src_sample_acks(0)  <= u64_true_divide_revised_CP_355_elements(126);
      u64_true_divide_revised_CP_355_elements(125)<= src_update_reqs(0);
      src_update_acks(0)  <= u64_true_divide_revised_CP_355_elements(127);
      u64_true_divide_revised_CP_355_elements(122) <= phi_mux_reqs(0);
      triggers(1)  <= u64_true_divide_revised_CP_355_elements(119);
      u64_true_divide_revised_CP_355_elements(128)<= src_sample_reqs(1);
      src_sample_acks(1)  <= u64_true_divide_revised_CP_355_elements(130);
      u64_true_divide_revised_CP_355_elements(129)<= src_update_reqs(1);
      src_update_acks(1)  <= u64_true_divide_revised_CP_355_elements(131);
      u64_true_divide_revised_CP_355_elements(120) <= phi_mux_reqs(1);
      phi_stmt_7532_phi_seq_706 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_7532_phi_seq_706") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => u64_true_divide_revised_CP_355_elements(115), 
          phi_sample_ack => u64_true_divide_revised_CP_355_elements(116), 
          phi_update_req => u64_true_divide_revised_CP_355_elements(117), 
          phi_update_ack => u64_true_divide_revised_CP_355_elements(118), 
          phi_mux_ack => u64_true_divide_revised_CP_355_elements(123), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_7536_phi_seq_760_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= u64_true_divide_revised_CP_355_elements(140);
      u64_true_divide_revised_CP_355_elements(143)<= src_sample_reqs(0);
      src_sample_acks(0)  <= u64_true_divide_revised_CP_355_elements(145);
      u64_true_divide_revised_CP_355_elements(144)<= src_update_reqs(0);
      src_update_acks(0)  <= u64_true_divide_revised_CP_355_elements(146);
      u64_true_divide_revised_CP_355_elements(141) <= phi_mux_reqs(0);
      triggers(1)  <= u64_true_divide_revised_CP_355_elements(138);
      u64_true_divide_revised_CP_355_elements(147)<= src_sample_reqs(1);
      src_sample_acks(1)  <= u64_true_divide_revised_CP_355_elements(149);
      u64_true_divide_revised_CP_355_elements(148)<= src_update_reqs(1);
      src_update_acks(1)  <= u64_true_divide_revised_CP_355_elements(150);
      u64_true_divide_revised_CP_355_elements(139) <= phi_mux_reqs(1);
      phi_stmt_7536_phi_seq_760 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_7536_phi_seq_760") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => u64_true_divide_revised_CP_355_elements(134), 
          phi_sample_ack => u64_true_divide_revised_CP_355_elements(135), 
          phi_update_req => u64_true_divide_revised_CP_355_elements(136), 
          phi_update_ack => u64_true_divide_revised_CP_355_elements(137), 
          phi_mux_ack => u64_true_divide_revised_CP_355_elements(142), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_397_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= u64_true_divide_revised_CP_355_elements(9);
        preds(1)  <= u64_true_divide_revised_CP_355_elements(10);
        entry_tmerge_397 : transition_merge -- 
          generic map(name => " entry_tmerge_397")
          port map (preds => preds, symbol_out => u64_true_divide_revised_CP_355_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u33_7493_wire : std_logic_vector(32 downto 0);
    signal CONCAT_u1_u65_7523_wire : std_logic_vector(64 downto 0);
    signal COUNT_7524 : std_logic_vector(7 downto 0);
    signal DIVIDEND_7518 : std_logic_vector(64 downto 0);
    signal INITIAL_QMASK_7489 : std_logic_vector(63 downto 0);
    signal INITIAL_QMASK_7489_7512_buffered : std_logic_vector(63 downto 0);
    signal NCOUNT_7555 : std_logic_vector(7 downto 0);
    signal NDIVIDEND_7555 : std_logic_vector(64 downto 0);
    signal NNCOUNT_7567 : std_logic_vector(7 downto 0);
    signal NNCOUNT_7567_7527_buffered : std_logic_vector(7 downto 0);
    signal NNDIVIDEND_7567 : std_logic_vector(64 downto 0);
    signal NNDIVIDEND_7567_7520_buffered : std_logic_vector(64 downto 0);
    signal NNQMASK_7567 : std_logic_vector(63 downto 0);
    signal NNQMASK_7567_7513_buffered : std_logic_vector(63 downto 0);
    signal NNQUOTIENT_7567 : std_logic_vector(63 downto 0);
    signal NNQUOTIENT_7567_7517_buffered : std_logic_vector(63 downto 0);
    signal NQMASK_7555 : std_logic_vector(63 downto 0);
    signal NQUOTIENT_7555 : std_logic_vector(63 downto 0);
    signal QMASK_7510 : std_logic_vector(63 downto 0);
    signal QUOTIENT_7514 : std_logic_vector(63 downto 0);
    signal R_ZERO_1_7491_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_7494_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_7521_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_2_7498_wire_constant : std_logic_vector(1 downto 0);
    signal R_ZERO_64_7516_wire_constant : std_logic_vector(63 downto 0);
    signal R_ZERO_8_7526_wire_constant : std_logic_vector(7 downto 0);
    signal SHIFTED_DIVIDEND_7489 : std_logic_vector(63 downto 0);
    signal SHIFTED_DIVISOR_34_2X_7501 : std_logic_vector(33 downto 0);
    signal SHIFTED_DIVISOR_34_2X_7501_7538_buffered : std_logic_vector(33 downto 0);
    signal SHIFTED_DIVISOR_34_2X_7501_7539_buffered : std_logic_vector(33 downto 0);
    signal SHIFTED_DIVISOR_34_3X_7506 : std_logic_vector(33 downto 0);
    signal SHIFTED_DIVISOR_34_3X_7506_7534_buffered : std_logic_vector(33 downto 0);
    signal SHIFTED_DIVISOR_34_3X_7506_7535_buffered : std_logic_vector(33 downto 0);
    signal SHIFTED_DIVISOR_34_7496 : std_logic_vector(33 downto 0);
    signal SHIFTED_DIVISOR_34_7496_7530_buffered : std_logic_vector(33 downto 0);
    signal SHIFTED_DIVISOR_34_7496_7531_buffered : std_logic_vector(33 downto 0);
    signal SHIFTED_DIVISOR_7489 : std_logic_vector(31 downto 0);
    signal U2X_7536 : std_logic_vector(33 downto 0);
    signal U3X_7532 : std_logic_vector(33 downto 0);
    signal U_7528 : std_logic_vector(33 downto 0);
    signal continue_flag_7572 : std_logic_vector(0 downto 0);
    signal konst_7570_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_ZERO_1_7491_wire_constant <= "0";
    R_ZERO_1_7494_wire_constant <= "0";
    R_ZERO_1_7521_wire_constant <= "0";
    R_ZERO_2_7498_wire_constant <= "00";
    R_ZERO_64_7516_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    R_ZERO_8_7526_wire_constant <= "00000000";
    konst_7570_wire_constant <= "00100001";
    phi_stmt_7510: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= INITIAL_QMASK_7489_7512_buffered & NNQMASK_7567_7513_buffered;
      req <= phi_stmt_7510_req_0 & phi_stmt_7510_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_7510",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_7510_ack_0,
          idata => idata,
          odata => QMASK_7510,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_7510
    phi_stmt_7514: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_64_7516_wire_constant & NNQUOTIENT_7567_7517_buffered;
      req <= phi_stmt_7514_req_0 & phi_stmt_7514_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_7514",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_7514_ack_0,
          idata => idata,
          odata => QUOTIENT_7514,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_7514
    phi_stmt_7518: Block -- phi operator 
      signal idata: std_logic_vector(129 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= NNDIVIDEND_7567_7520_buffered & CONCAT_u1_u65_7523_wire;
      req <= phi_stmt_7518_req_0 & phi_stmt_7518_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_7518",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 65) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_7518_ack_0,
          idata => idata,
          odata => DIVIDEND_7518,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_7518
    phi_stmt_7524: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_7526_wire_constant & NNCOUNT_7567_7527_buffered;
      req <= phi_stmt_7524_req_0 & phi_stmt_7524_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_7524",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_7524_ack_0,
          idata => idata,
          odata => COUNT_7524,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_7524
    phi_stmt_7528: Block -- phi operator 
      signal idata: std_logic_vector(67 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= SHIFTED_DIVISOR_34_7496_7530_buffered & SHIFTED_DIVISOR_34_7496_7531_buffered;
      req <= phi_stmt_7528_req_0 & phi_stmt_7528_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_7528",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 34) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_7528_ack_0,
          idata => idata,
          odata => U_7528,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_7528
    phi_stmt_7532: Block -- phi operator 
      signal idata: std_logic_vector(67 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= SHIFTED_DIVISOR_34_3X_7506_7534_buffered & SHIFTED_DIVISOR_34_3X_7506_7535_buffered;
      req <= phi_stmt_7532_req_0 & phi_stmt_7532_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_7532",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 34) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_7532_ack_0,
          idata => idata,
          odata => U3X_7532,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_7532
    phi_stmt_7536: Block -- phi operator 
      signal idata: std_logic_vector(67 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= SHIFTED_DIVISOR_34_2X_7501_7538_buffered & SHIFTED_DIVISOR_34_2X_7501_7539_buffered;
      req <= phi_stmt_7536_req_0 & phi_stmt_7536_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_7536",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 34) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_7536_ack_0,
          idata => idata,
          odata => U2X_7536,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_7536
    INITIAL_QMASK_7489_7512_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= INITIAL_QMASK_7489_7512_buf_req_0;
      INITIAL_QMASK_7489_7512_buf_ack_0<= wack(0);
      rreq(0) <= INITIAL_QMASK_7489_7512_buf_req_1;
      INITIAL_QMASK_7489_7512_buf_ack_1<= rack(0);
      INITIAL_QMASK_7489_7512_buf : InterlockBuffer generic map ( -- 
        name => "INITIAL_QMASK_7489_7512_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => INITIAL_QMASK_7489,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => INITIAL_QMASK_7489_7512_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    NNCOUNT_7567_7527_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NNCOUNT_7567_7527_buf_req_0;
      NNCOUNT_7567_7527_buf_ack_0<= wack(0);
      rreq(0) <= NNCOUNT_7567_7527_buf_req_1;
      NNCOUNT_7567_7527_buf_ack_1<= rack(0);
      NNCOUNT_7567_7527_buf : InterlockBuffer generic map ( -- 
        name => "NNCOUNT_7567_7527_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NNCOUNT_7567,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NNCOUNT_7567_7527_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    NNDIVIDEND_7567_7520_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NNDIVIDEND_7567_7520_buf_req_0;
      NNDIVIDEND_7567_7520_buf_ack_0<= wack(0);
      rreq(0) <= NNDIVIDEND_7567_7520_buf_req_1;
      NNDIVIDEND_7567_7520_buf_ack_1<= rack(0);
      NNDIVIDEND_7567_7520_buf : InterlockBuffer generic map ( -- 
        name => "NNDIVIDEND_7567_7520_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 65,
        out_data_width => 65,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NNDIVIDEND_7567,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NNDIVIDEND_7567_7520_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    NNQMASK_7567_7513_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NNQMASK_7567_7513_buf_req_0;
      NNQMASK_7567_7513_buf_ack_0<= wack(0);
      rreq(0) <= NNQMASK_7567_7513_buf_req_1;
      NNQMASK_7567_7513_buf_ack_1<= rack(0);
      NNQMASK_7567_7513_buf : InterlockBuffer generic map ( -- 
        name => "NNQMASK_7567_7513_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NNQMASK_7567,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NNQMASK_7567_7513_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    NNQUOTIENT_7567_7517_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NNQUOTIENT_7567_7517_buf_req_0;
      NNQUOTIENT_7567_7517_buf_ack_0<= wack(0);
      rreq(0) <= NNQUOTIENT_7567_7517_buf_req_1;
      NNQUOTIENT_7567_7517_buf_ack_1<= rack(0);
      NNQUOTIENT_7567_7517_buf : InterlockBuffer generic map ( -- 
        name => "NNQUOTIENT_7567_7517_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NNQUOTIENT_7567,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NNQUOTIENT_7567_7517_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    SHIFTED_DIVISOR_34_2X_7501_7538_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= SHIFTED_DIVISOR_34_2X_7501_7538_buf_req_0;
      SHIFTED_DIVISOR_34_2X_7501_7538_buf_ack_0<= wack(0);
      rreq(0) <= SHIFTED_DIVISOR_34_2X_7501_7538_buf_req_1;
      SHIFTED_DIVISOR_34_2X_7501_7538_buf_ack_1<= rack(0);
      SHIFTED_DIVISOR_34_2X_7501_7538_buf : InterlockBuffer generic map ( -- 
        name => "SHIFTED_DIVISOR_34_2X_7501_7538_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 34,
        out_data_width => 34,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => SHIFTED_DIVISOR_34_2X_7501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => SHIFTED_DIVISOR_34_2X_7501_7538_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    SHIFTED_DIVISOR_34_2X_7501_7539_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= SHIFTED_DIVISOR_34_2X_7501_7539_buf_req_0;
      SHIFTED_DIVISOR_34_2X_7501_7539_buf_ack_0<= wack(0);
      rreq(0) <= SHIFTED_DIVISOR_34_2X_7501_7539_buf_req_1;
      SHIFTED_DIVISOR_34_2X_7501_7539_buf_ack_1<= rack(0);
      SHIFTED_DIVISOR_34_2X_7501_7539_buf : InterlockBuffer generic map ( -- 
        name => "SHIFTED_DIVISOR_34_2X_7501_7539_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 34,
        out_data_width => 34,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => SHIFTED_DIVISOR_34_2X_7501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => SHIFTED_DIVISOR_34_2X_7501_7539_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    SHIFTED_DIVISOR_34_3X_7506_7534_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= SHIFTED_DIVISOR_34_3X_7506_7534_buf_req_0;
      SHIFTED_DIVISOR_34_3X_7506_7534_buf_ack_0<= wack(0);
      rreq(0) <= SHIFTED_DIVISOR_34_3X_7506_7534_buf_req_1;
      SHIFTED_DIVISOR_34_3X_7506_7534_buf_ack_1<= rack(0);
      SHIFTED_DIVISOR_34_3X_7506_7534_buf : InterlockBuffer generic map ( -- 
        name => "SHIFTED_DIVISOR_34_3X_7506_7534_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 34,
        out_data_width => 34,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => SHIFTED_DIVISOR_34_3X_7506,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => SHIFTED_DIVISOR_34_3X_7506_7534_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    SHIFTED_DIVISOR_34_3X_7506_7535_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= SHIFTED_DIVISOR_34_3X_7506_7535_buf_req_0;
      SHIFTED_DIVISOR_34_3X_7506_7535_buf_ack_0<= wack(0);
      rreq(0) <= SHIFTED_DIVISOR_34_3X_7506_7535_buf_req_1;
      SHIFTED_DIVISOR_34_3X_7506_7535_buf_ack_1<= rack(0);
      SHIFTED_DIVISOR_34_3X_7506_7535_buf : InterlockBuffer generic map ( -- 
        name => "SHIFTED_DIVISOR_34_3X_7506_7535_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 34,
        out_data_width => 34,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => SHIFTED_DIVISOR_34_3X_7506,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => SHIFTED_DIVISOR_34_3X_7506_7535_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    SHIFTED_DIVISOR_34_7496_7530_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= SHIFTED_DIVISOR_34_7496_7530_buf_req_0;
      SHIFTED_DIVISOR_34_7496_7530_buf_ack_0<= wack(0);
      rreq(0) <= SHIFTED_DIVISOR_34_7496_7530_buf_req_1;
      SHIFTED_DIVISOR_34_7496_7530_buf_ack_1<= rack(0);
      SHIFTED_DIVISOR_34_7496_7530_buf : InterlockBuffer generic map ( -- 
        name => "SHIFTED_DIVISOR_34_7496_7530_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 34,
        out_data_width => 34,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => SHIFTED_DIVISOR_34_7496,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => SHIFTED_DIVISOR_34_7496_7530_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    SHIFTED_DIVISOR_34_7496_7531_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= SHIFTED_DIVISOR_34_7496_7531_buf_req_0;
      SHIFTED_DIVISOR_34_7496_7531_buf_ack_0<= wack(0);
      rreq(0) <= SHIFTED_DIVISOR_34_7496_7531_buf_req_1;
      SHIFTED_DIVISOR_34_7496_7531_buf_ack_1<= rack(0);
      SHIFTED_DIVISOR_34_7496_7531_buf : InterlockBuffer generic map ( -- 
        name => "SHIFTED_DIVISOR_34_7496_7531_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 34,
        out_data_width => 34,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => SHIFTED_DIVISOR_34_7496,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => SHIFTED_DIVISOR_34_7496_7531_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_quotient_7576_inst
    process(NNQUOTIENT_7567) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := NNQUOTIENT_7567(63 downto 0);
      quotient_buffer <= tmp_var; -- 
    end process;
    do_while_stmt_7508_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_7572;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_7508_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_7508_branch_req_0,
          ack0 => do_while_stmt_7508_branch_ack_0,
          ack1 => do_while_stmt_7508_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator ADD_u34_u34_7505_inst
    SHIFTED_DIVISOR_34_3X_7506 <= std_logic_vector(unsigned(SHIFTED_DIVISOR_34_7496) + unsigned(SHIFTED_DIVISOR_34_2X_7501));
    -- flow through binary operator CONCAT_u1_u33_7493_inst
    process(R_ZERO_1_7491_wire_constant, SHIFTED_DIVISOR_7489) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_1_7491_wire_constant, SHIFTED_DIVISOR_7489, tmp_var);
      CONCAT_u1_u33_7493_wire <= tmp_var; --
    end process;
    -- shared split operator group (2) : CONCAT_u1_u65_7523_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(64 downto 0);
      signal data_out: std_logic_vector(64 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ZERO_1_7521_wire_constant & SHIFTED_DIVIDEND_7489;
      CONCAT_u1_u65_7523_wire <= data_out(64 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u1_u65_7523_inst_req_0;
      CONCAT_u1_u65_7523_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u1_u65_7523_inst_req_1;
      CONCAT_u1_u65_7523_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_2_gI: SplitGuardInterface generic map(name => "ApConcat_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 65,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- flow through binary operator CONCAT_u2_u34_7500_inst
    process(R_ZERO_2_7498_wire_constant, SHIFTED_DIVISOR_7489) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_2_7498_wire_constant, SHIFTED_DIVISOR_7489, tmp_var);
      SHIFTED_DIVISOR_34_2X_7501 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u33_u34_7495_inst
    process(CONCAT_u1_u33_7493_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u33_7493_wire, R_ZERO_1_7494_wire_constant, tmp_var);
      SHIFTED_DIVISOR_34_7496 <= tmp_var; --
    end process;
    -- flow through binary operator ULT_u8_u1_7571_inst
    process(NNCOUNT_7567) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(NNCOUNT_7567, konst_7570_wire_constant, tmp_var);
      continue_flag_7572 <= tmp_var; --
    end process;
    operator_alignDivisorToDividendRevised_6697_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_7489_call_req_0;
      call_stmt_7489_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_7489_call_req_1;
      call_stmt_7489_call_ack_1<= update_ack(0);
      call_stmt_7489_call: alignDivisorToDividendRevised_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        DIVIDEND => udividend_buffer,
        udivisor => udivisor_buffer,
        SHIFTED_DIVIDEND => SHIFTED_DIVIDEND_7489,
        SHIFTED_DIVISOR => SHIFTED_DIVISOR_7489,
        INITIAL_QMASK => INITIAL_QMASK_7489,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    volatile_operator_u64_true_divide_revised_core_6722: u64_true_divide_revised_core_Volatile port map(QMASK => QMASK_7510, QUOTIENT => QUOTIENT_7514, DIVIDEND => DIVIDEND_7518, SHIFTED_DIVISOR_34 => U_7528, SHIFTED_DIVISOR_34_2X => U2X_7536, SHIFTED_DIVISOR_34_3X => U3X_7532, COUNT => COUNT_7524, NQMASK => NQMASK_7555, NQUOTIENT => NQUOTIENT_7555, NDIVIDEND => NDIVIDEND_7555, NCOUNT => NCOUNT_7555); 
    volatile_operator_u64_true_divide_revised_core_6723: u64_true_divide_revised_core_Volatile port map(QMASK => NQMASK_7555, QUOTIENT => NQUOTIENT_7555, DIVIDEND => NDIVIDEND_7555, SHIFTED_DIVISOR_34 => U_7528, SHIFTED_DIVISOR_34_2X => U2X_7536, SHIFTED_DIVISOR_34_3X => U3X_7532, COUNT => NCOUNT_7555, NQMASK => NNQMASK_7567, NQUOTIENT => NNQUOTIENT_7567, NDIVIDEND => NNDIVIDEND_7567, NCOUNT => NNCOUNT_7567); 
    -- 
  end Block; -- data_path
  -- 
end u64_true_divide_revised_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity u64_true_divide_revised_core_Volatile is -- 
  port ( -- 
    QMASK : in  std_logic_vector(63 downto 0);
    QUOTIENT : in  std_logic_vector(63 downto 0);
    DIVIDEND : in  std_logic_vector(64 downto 0);
    SHIFTED_DIVISOR_34 : in  std_logic_vector(33 downto 0);
    SHIFTED_DIVISOR_34_2X : in  std_logic_vector(33 downto 0);
    SHIFTED_DIVISOR_34_3X : in  std_logic_vector(33 downto 0);
    COUNT : in  std_logic_vector(7 downto 0);
    NQMASK : out  std_logic_vector(63 downto 0);
    NQUOTIENT : out  std_logic_vector(63 downto 0);
    NDIVIDEND : out  std_logic_vector(64 downto 0);
    NCOUNT : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity u64_true_divide_revised_core_Volatile;
architecture u64_true_divide_revised_core_Volatile_arch of u64_true_divide_revised_core_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(303-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal QMASK_buffer :  std_logic_vector(63 downto 0);
  signal QUOTIENT_buffer :  std_logic_vector(63 downto 0);
  signal DIVIDEND_buffer :  std_logic_vector(64 downto 0);
  signal SHIFTED_DIVISOR_34_buffer :  std_logic_vector(33 downto 0);
  signal SHIFTED_DIVISOR_34_2X_buffer :  std_logic_vector(33 downto 0);
  signal SHIFTED_DIVISOR_34_3X_buffer :  std_logic_vector(33 downto 0);
  signal COUNT_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal NQMASK_buffer :  std_logic_vector(63 downto 0);
  signal NQUOTIENT_buffer :  std_logic_vector(63 downto 0);
  signal NDIVIDEND_buffer :  std_logic_vector(64 downto 0);
  signal NCOUNT_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  component u_cmp_34_Volatile is -- 
    port ( -- 
      a : in  std_logic_vector(33 downto 0);
      b : in  std_logic_vector(33 downto 0);
      l : out  std_logic_vector(0 downto 0);
      g : out  std_logic_vector(0 downto 0);
      e : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  QMASK_buffer <= QMASK;
  QUOTIENT_buffer <= QUOTIENT;
  DIVIDEND_buffer <= DIVIDEND;
  SHIFTED_DIVISOR_34_buffer <= SHIFTED_DIVISOR_34;
  SHIFTED_DIVISOR_34_2X_buffer <= SHIFTED_DIVISOR_34_2X;
  SHIFTED_DIVISOR_34_3X_buffer <= SHIFTED_DIVISOR_34_3X;
  COUNT_buffer <= COUNT;
  -- output handling  -------------------------------------------------------
  NQMASK <= NQMASK_buffer;
  NQUOTIENT <= NQUOTIENT_buffer;
  NDIVIDEND <= NDIVIDEND_buffer;
  NCOUNT <= NCOUNT_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal MUX_7440_wire : std_logic_vector(33 downto 0);
    signal MUX_7441_wire : std_logic_vector(33 downto 0);
    signal MUX_7454_wire : std_logic_vector(63 downto 0);
    signal MUX_7455_wire : std_logic_vector(63 downto 0);
    signal OR_u64_u64_7448_wire : std_logic_vector(63 downto 0);
    signal QMASK_RS_1_7384 : std_logic_vector(63 downto 0);
    signal QMASK_RS_2_7390 : std_logic_vector(63 downto 0);
    signal R_ZERO_1_7380_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_1_7386_wire_constant : std_logic_vector(0 downto 0);
    signal R_ZERO_2_7473_wire_constant : std_logic_vector(1 downto 0);
    signal SUB_u34_u34_7461_wire : std_logic_vector(33 downto 0);
    signal div_h_34_7394 : std_logic_vector(33 downto 0);
    signal div_l_31_7398 : std_logic_vector(30 downto 0);
    signal dividend_minus_divisor_7464 : std_logic_vector(64 downto 0);
    signal e_2x_7410 : std_logic_vector(0 downto 0);
    signal e_3x_7416 : std_logic_vector(0 downto 0);
    signal e_x_7404 : std_logic_vector(0 downto 0);
    signal g_2x_7410 : std_logic_vector(0 downto 0);
    signal g_3x_7416 : std_logic_vector(0 downto 0);
    signal g_x_7404 : std_logic_vector(0 downto 0);
    signal ge_2X_7426 : std_logic_vector(0 downto 0);
    signal ge_3X_7431 : std_logic_vector(0 downto 0);
    signal ge_X_7421 : std_logic_vector(0 downto 0);
    signal konst_7376_wire_constant : std_logic_vector(7 downto 0);
    signal konst_7439_wire_constant : std_logic_vector(33 downto 0);
    signal konst_7453_wire_constant : std_logic_vector(63 downto 0);
    signal l_2x_7410 : std_logic_vector(0 downto 0);
    signal l_3x_7416 : std_logic_vector(0 downto 0);
    signal l_x_7404 : std_logic_vector(0 downto 0);
    signal qmask_val_7457 : std_logic_vector(63 downto 0);
    signal slice_7382_wire : std_logic_vector(62 downto 0);
    signal slice_7388_wire : std_logic_vector(62 downto 0);
    signal slice_7472_wire : std_logic_vector(62 downto 0);
    signal sub_val_7443 : std_logic_vector(33 downto 0);
    -- 
  begin -- 
    R_ZERO_1_7380_wire_constant <= "0";
    R_ZERO_1_7386_wire_constant <= "0";
    R_ZERO_2_7473_wire_constant <= "00";
    konst_7376_wire_constant <= "00000010";
    konst_7439_wire_constant <= "0000000000000000000000000000000000";
    konst_7453_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- flow-through select operator MUX_7440_inst
    MUX_7440_wire <= SHIFTED_DIVISOR_34_2X_buffer when (ge_2X_7426(0) /=  '0') else konst_7439_wire_constant;
    -- flow-through select operator MUX_7441_inst
    MUX_7441_wire <= SHIFTED_DIVISOR_34_buffer when (ge_X_7421(0) /=  '0') else MUX_7440_wire;
    -- flow-through select operator MUX_7442_inst
    sub_val_7443 <= SHIFTED_DIVISOR_34_3X_buffer when (ge_3X_7431(0) /=  '0') else MUX_7441_wire;
    -- flow-through select operator MUX_7454_inst
    MUX_7454_wire <= QMASK_RS_1_7384 when (ge_2X_7426(0) /=  '0') else konst_7453_wire_constant;
    -- flow-through select operator MUX_7455_inst
    MUX_7455_wire <= QMASK_buffer when (ge_X_7421(0) /=  '0') else MUX_7454_wire;
    -- flow-through select operator MUX_7456_inst
    qmask_val_7457 <= OR_u64_u64_7448_wire when (ge_3X_7431(0) /=  '0') else MUX_7455_wire;
    -- flow-through slice operator slice_7382_inst
    slice_7382_wire <= QMASK_buffer(63 downto 1);
    -- flow-through slice operator slice_7388_inst
    slice_7388_wire <= QMASK_RS_1_7384(63 downto 1);
    -- flow-through slice operator slice_7393_inst
    div_h_34_7394 <= DIVIDEND_buffer(64 downto 31);
    -- flow-through slice operator slice_7397_inst
    div_l_31_7398 <= DIVIDEND_buffer(30 downto 0);
    -- flow-through slice operator slice_7472_inst
    slice_7472_wire <= dividend_minus_divisor_7464(62 downto 0);
    -- interlock W_NQMASK_7476_inst
    process(QMASK_RS_2_7390) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := QMASK_RS_2_7390(63 downto 0);
      NQMASK_buffer <= tmp_var; -- 
    end process;
    -- flow through binary operator ADD_u8_u8_7377_inst
    NCOUNT_buffer <= std_logic_vector(unsigned(COUNT_buffer) + unsigned(konst_7376_wire_constant));
    -- flow through binary operator CONCAT_u1_u64_7383_inst
    process(R_ZERO_1_7380_wire_constant, slice_7382_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_1_7380_wire_constant, slice_7382_wire, tmp_var);
      QMASK_RS_1_7384 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u64_7389_inst
    process(R_ZERO_1_7386_wire_constant, slice_7388_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ZERO_1_7386_wire_constant, slice_7388_wire, tmp_var);
      QMASK_RS_2_7390 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u34_u65_7463_inst
    process(SUB_u34_u34_7461_wire, div_l_31_7398) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(SUB_u34_u34_7461_wire, div_l_31_7398, tmp_var);
      dividend_minus_divisor_7464 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u63_u65_7474_inst
    process(slice_7472_wire) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_7472_wire, R_ZERO_2_7473_wire_constant, tmp_var);
      NDIVIDEND_buffer <= tmp_var; --
    end process;
    -- flow through binary operator OR_u1_u1_7420_inst
    ge_X_7421 <= (g_x_7404 or e_x_7404);
    -- flow through binary operator OR_u1_u1_7425_inst
    ge_2X_7426 <= (g_2x_7410 or e_2x_7410);
    -- flow through binary operator OR_u1_u1_7430_inst
    ge_3X_7431 <= (g_3x_7416 or e_3x_7416);
    -- flow through binary operator OR_u64_u64_7448_inst
    OR_u64_u64_7448_wire <= (QMASK_buffer or QMASK_RS_1_7384);
    -- flow through binary operator OR_u64_u64_7468_inst
    NQUOTIENT_buffer <= (QUOTIENT_buffer or qmask_val_7457);
    -- flow through binary operator SUB_u34_u34_7461_inst
    SUB_u34_u34_7461_wire <= std_logic_vector(unsigned(div_h_34_7394) - unsigned(sub_val_7443));
    volatile_operator_u_cmp_34_6205: u_cmp_34_Volatile port map(a => div_h_34_7394, b => SHIFTED_DIVISOR_34_buffer, l => l_x_7404, g => g_x_7404, e => e_x_7404); 
    volatile_operator_u_cmp_34_6206: u_cmp_34_Volatile port map(a => div_h_34_7394, b => SHIFTED_DIVISOR_34_2X_buffer, l => l_2x_7410, g => g_2x_7410, e => e_2x_7410); 
    volatile_operator_u_cmp_34_6207: u_cmp_34_Volatile port map(a => div_h_34_7394, b => SHIFTED_DIVISOR_34_3X_buffer, l => l_3x_7416, g => g_3x_7416, e => e_3x_7416); 
    -- 
  end Block; -- data_path
  -- 
end u64_true_divide_revised_core_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity u_cmp_32_Volatile is -- 
  port ( -- 
    a : in  std_logic_vector(31 downto 0);
    b : in  std_logic_vector(31 downto 0);
    l : out  std_logic_vector(0 downto 0);
    g : out  std_logic_vector(0 downto 0);
    e : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity u_cmp_32_Volatile;
architecture u_cmp_32_Volatile_arch of u_cmp_32_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(64-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal a_buffer :  std_logic_vector(31 downto 0);
  signal b_buffer :  std_logic_vector(31 downto 0);
  -- output port buffer signals
  signal l_buffer :  std_logic_vector(0 downto 0);
  signal g_buffer :  std_logic_vector(0 downto 0);
  signal e_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  a_buffer <= a;
  b_buffer <= b;
  -- output handling  -------------------------------------------------------
  l <= l_buffer;
  g <= g_buffer;
  e <= e_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1254_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1266_wire : std_logic_vector(0 downto 0);
    signal ah_1211 : std_logic_vector(15 downto 0);
    signal al_1207 : std_logic_vector(15 downto 0);
    signal bh_1219 : std_logic_vector(15 downto 0);
    signal bl_1215 : std_logic_vector(15 downto 0);
    signal eh_1249 : std_logic_vector(0 downto 0);
    signal el_1234 : std_logic_vector(0 downto 0);
    signal gh_1244 : std_logic_vector(0 downto 0);
    signal gl_1229 : std_logic_vector(0 downto 0);
    signal lh_1239 : std_logic_vector(0 downto 0);
    signal ll_1224 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_1206_inst
    al_1207 <= a_buffer(15 downto 0);
    -- flow-through slice operator slice_1210_inst
    ah_1211 <= a_buffer(31 downto 16);
    -- flow-through slice operator slice_1214_inst
    bl_1215 <= b_buffer(15 downto 0);
    -- flow-through slice operator slice_1218_inst
    bh_1219 <= b_buffer(31 downto 16);
    -- flow through binary operator AND_u1_u1_1254_inst
    AND_u1_u1_1254_wire <= (eh_1249 and ll_1224);
    -- flow through binary operator AND_u1_u1_1260_inst
    e_buffer <= (eh_1249 and el_1234);
    -- flow through binary operator AND_u1_u1_1266_inst
    AND_u1_u1_1266_wire <= (eh_1249 and gl_1229);
    -- flow through binary operator EQ_u16_u1_1233_inst
    process(al_1207, bl_1215) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(al_1207, bl_1215, tmp_var);
      el_1234 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u16_u1_1248_inst
    process(ah_1211, bh_1219) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ah_1211, bh_1219, tmp_var);
      eh_1249 <= tmp_var; --
    end process;
    -- flow through binary operator OR_u1_u1_1255_inst
    l_buffer <= (lh_1239 or AND_u1_u1_1254_wire);
    -- flow through binary operator OR_u1_u1_1267_inst
    g_buffer <= (gh_1244 or AND_u1_u1_1266_wire);
    -- flow through binary operator UGT_u16_u1_1228_inst
    process(al_1207, bl_1215) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(al_1207, bl_1215, tmp_var);
      gl_1229 <= tmp_var; --
    end process;
    -- flow through binary operator UGT_u16_u1_1243_inst
    process(ah_1211, bh_1219) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ah_1211, bh_1219, tmp_var);
      gh_1244 <= tmp_var; --
    end process;
    -- flow through binary operator ULT_u16_u1_1223_inst
    process(al_1207, bl_1215) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(al_1207, bl_1215, tmp_var);
      ll_1224 <= tmp_var; --
    end process;
    -- flow through binary operator ULT_u16_u1_1238_inst
    process(ah_1211, bh_1219) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(ah_1211, bh_1219, tmp_var);
      lh_1239 <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end u_cmp_32_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity u_cmp_34_Volatile is -- 
  port ( -- 
    a : in  std_logic_vector(33 downto 0);
    b : in  std_logic_vector(33 downto 0);
    l : out  std_logic_vector(0 downto 0);
    g : out  std_logic_vector(0 downto 0);
    e : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity u_cmp_34_Volatile;
architecture u_cmp_34_Volatile_arch of u_cmp_34_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(68-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal a_buffer :  std_logic_vector(33 downto 0);
  signal b_buffer :  std_logic_vector(33 downto 0);
  -- output port buffer signals
  signal l_buffer :  std_logic_vector(0 downto 0);
  signal g_buffer :  std_logic_vector(0 downto 0);
  signal e_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  component u_cmp_32_Volatile is -- 
    port ( -- 
      a : in  std_logic_vector(31 downto 0);
      b : in  std_logic_vector(31 downto 0);
      l : out  std_logic_vector(0 downto 0);
      g : out  std_logic_vector(0 downto 0);
      e : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  a_buffer <= a;
  b_buffer <= b;
  -- output handling  -------------------------------------------------------
  l <= l_buffer;
  g <= g_buffer;
  e <= e_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_7345_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_7357_wire : std_logic_vector(0 downto 0);
    signal ah_7311 : std_logic_vector(1 downto 0);
    signal al_7307 : std_logic_vector(31 downto 0);
    signal bh_7319 : std_logic_vector(1 downto 0);
    signal bl_7315 : std_logic_vector(31 downto 0);
    signal eh_7340 : std_logic_vector(0 downto 0);
    signal el_7325 : std_logic_vector(0 downto 0);
    signal gh_7335 : std_logic_vector(0 downto 0);
    signal gl_7325 : std_logic_vector(0 downto 0);
    signal lh_7330 : std_logic_vector(0 downto 0);
    signal ll_7325 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_7306_inst
    al_7307 <= a_buffer(31 downto 0);
    -- flow-through slice operator slice_7310_inst
    ah_7311 <= a_buffer(33 downto 32);
    -- flow-through slice operator slice_7314_inst
    bl_7315 <= b_buffer(31 downto 0);
    -- flow-through slice operator slice_7318_inst
    bh_7319 <= b_buffer(33 downto 32);
    -- flow through binary operator AND_u1_u1_7345_inst
    AND_u1_u1_7345_wire <= (eh_7340 and ll_7325);
    -- flow through binary operator AND_u1_u1_7351_inst
    e_buffer <= (eh_7340 and el_7325);
    -- flow through binary operator AND_u1_u1_7357_inst
    AND_u1_u1_7357_wire <= (eh_7340 and gl_7325);
    -- flow through binary operator EQ_u2_u1_7339_inst
    process(ah_7311, bh_7319) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ah_7311, bh_7319, tmp_var);
      eh_7340 <= tmp_var; --
    end process;
    -- flow through binary operator OR_u1_u1_7346_inst
    l_buffer <= (lh_7330 or AND_u1_u1_7345_wire);
    -- flow through binary operator OR_u1_u1_7358_inst
    g_buffer <= (gh_7335 or AND_u1_u1_7357_wire);
    -- flow through binary operator UGT_u2_u1_7334_inst
    process(ah_7311, bh_7319) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ah_7311, bh_7319, tmp_var);
      gh_7335 <= tmp_var; --
    end process;
    -- flow through binary operator ULT_u2_u1_7329_inst
    process(ah_7311, bh_7319) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(ah_7311, bh_7319, tmp_var);
      lh_7330 <= tmp_var; --
    end process;
    volatile_operator_u_cmp_32_6132: u_cmp_32_Volatile port map(a => al_7307, b => bl_7315, l => ll_7325, g => gl_7325, e => el_7325); 
    -- 
  end Block; -- data_path
  -- 
end u_cmp_34_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity u_set_index_64_Volatile is -- 
  port ( -- 
    idx : in  std_logic_vector(5 downto 0);
    x : out  std_logic_vector(63 downto 0)-- 
  );
  -- 
end entity u_set_index_64_Volatile;
architecture u_set_index_64_Volatile_arch of u_set_index_64_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(6-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal idx_buffer :  std_logic_vector(5 downto 0);
  -- output port buffer signals
  signal x_buffer :  std_logic_vector(63 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  idx_buffer <= idx;
  -- output handling  -------------------------------------------------------
  x <= x_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u16_u32_1379_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1382_wire : std_logic_vector(31 downto 0);
    signal R_ZERO_16_1347_wire_constant : std_logic_vector(15 downto 0);
    signal R_ZERO_16_1360_wire_constant : std_logic_vector(15 downto 0);
    signal R_ZERO_16_1373_wire_constant : std_logic_vector(15 downto 0);
    signal SHL_u16_u16_1346_wire : std_logic_vector(15 downto 0);
    signal SHL_u16_u16_1359_wire : std_logic_vector(15 downto 0);
    signal SHL_u16_u16_1372_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_1345_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_1358_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_1371_wire : std_logic_vector(15 downto 0);
    signal UGE_u16_u1_1340_wire : std_logic_vector(0 downto 0);
    signal UGE_u16_u1_1353_wire : std_logic_vector(0 downto 0);
    signal UGE_u16_u1_1366_wire : std_logic_vector(0 downto 0);
    signal idx_16_1330 : std_logic_vector(15 downto 0);
    signal konst_1339_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1344_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1352_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1357_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1365_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1370_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1333_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1342_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1355_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1368_wire_constant : std_logic_vector(15 downto 0);
    signal x00_1336 : std_logic_vector(15 downto 0);
    signal x01_1349 : std_logic_vector(15 downto 0);
    signal x10_1362 : std_logic_vector(15 downto 0);
    signal x11_1375 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ZERO_16_1347_wire_constant <= "0000000000000000";
    R_ZERO_16_1360_wire_constant <= "0000000000000000";
    R_ZERO_16_1373_wire_constant <= "0000000000000000";
    konst_1339_wire_constant <= "0000000000010000";
    konst_1344_wire_constant <= "0000000000010000";
    konst_1352_wire_constant <= "0000000000100000";
    konst_1357_wire_constant <= "0000000000100000";
    konst_1365_wire_constant <= "0000000000110000";
    konst_1370_wire_constant <= "0000000000110000";
    type_cast_1333_wire_constant <= "0000000000000001";
    type_cast_1342_wire_constant <= "0000000000000001";
    type_cast_1355_wire_constant <= "0000000000000001";
    type_cast_1368_wire_constant <= "0000000000000001";
    -- flow-through select operator MUX_1348_inst
    x01_1349 <= SHL_u16_u16_1346_wire when (UGE_u16_u1_1340_wire(0) /=  '0') else R_ZERO_16_1347_wire_constant;
    -- flow-through select operator MUX_1361_inst
    x10_1362 <= SHL_u16_u16_1359_wire when (UGE_u16_u1_1353_wire(0) /=  '0') else R_ZERO_16_1360_wire_constant;
    -- flow-through select operator MUX_1374_inst
    x11_1375 <= SHL_u16_u16_1372_wire when (UGE_u16_u1_1366_wire(0) /=  '0') else R_ZERO_16_1373_wire_constant;
    -- interlock type_cast_1329_inst
    process(idx_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := idx_buffer(5 downto 0);
      idx_16_1330 <= tmp_var; -- 
    end process;
    -- flow through binary operator CONCAT_u16_u32_1379_inst
    process(x11_1375, x10_1362) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(x11_1375, x10_1362, tmp_var);
      CONCAT_u16_u32_1379_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u16_u32_1382_inst
    process(x01_1349, x00_1336) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(x01_1349, x00_1336, tmp_var);
      CONCAT_u16_u32_1382_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u32_u64_1383_inst
    process(CONCAT_u16_u32_1379_wire, CONCAT_u16_u32_1382_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u16_u32_1379_wire, CONCAT_u16_u32_1382_wire, tmp_var);
      x_buffer <= tmp_var; --
    end process;
    -- flow through binary operator SHL_u16_u16_1335_inst
    process(type_cast_1333_wire_constant, idx_16_1330) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(type_cast_1333_wire_constant, idx_16_1330, tmp_var);
      x00_1336 <= tmp_var; --
    end process;
    -- flow through binary operator SHL_u16_u16_1346_inst
    process(type_cast_1342_wire_constant, SUB_u16_u16_1345_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(type_cast_1342_wire_constant, SUB_u16_u16_1345_wire, tmp_var);
      SHL_u16_u16_1346_wire <= tmp_var; --
    end process;
    -- flow through binary operator SHL_u16_u16_1359_inst
    process(type_cast_1355_wire_constant, SUB_u16_u16_1358_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(type_cast_1355_wire_constant, SUB_u16_u16_1358_wire, tmp_var);
      SHL_u16_u16_1359_wire <= tmp_var; --
    end process;
    -- flow through binary operator SHL_u16_u16_1372_inst
    process(type_cast_1368_wire_constant, SUB_u16_u16_1371_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(type_cast_1368_wire_constant, SUB_u16_u16_1371_wire, tmp_var);
      SHL_u16_u16_1372_wire <= tmp_var; --
    end process;
    -- flow through binary operator SUB_u16_u16_1345_inst
    SUB_u16_u16_1345_wire <= std_logic_vector(unsigned(idx_16_1330) - unsigned(konst_1344_wire_constant));
    -- flow through binary operator SUB_u16_u16_1358_inst
    SUB_u16_u16_1358_wire <= std_logic_vector(unsigned(idx_16_1330) - unsigned(konst_1357_wire_constant));
    -- flow through binary operator SUB_u16_u16_1371_inst
    SUB_u16_u16_1371_wire <= std_logic_vector(unsigned(idx_16_1330) - unsigned(konst_1370_wire_constant));
    -- flow through binary operator UGE_u16_u1_1340_inst
    process(idx_16_1330) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(idx_16_1330, konst_1339_wire_constant, tmp_var);
      UGE_u16_u1_1340_wire <= tmp_var; --
    end process;
    -- flow through binary operator UGE_u16_u1_1353_inst
    process(idx_16_1330) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(idx_16_1330, konst_1352_wire_constant, tmp_var);
      UGE_u16_u1_1353_wire <= tmp_var; --
    end process;
    -- flow through binary operator UGE_u16_u1_1366_inst
    process(idx_16_1330) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(idx_16_1330, konst_1365_wire_constant, tmp_var);
      UGE_u16_u1_1366_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end u_set_index_64_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library iunit_exec;
use iunit_exec.iu_exec_global_package.all;
entity iu_exec is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    iunit_exec_fast_alu_result_to_writeback_pipe_read_data: out std_logic_vector(108 downto 0);
    iunit_exec_fast_alu_result_to_writeback_pipe_read_req : in std_logic_vector(0 downto 0);
    iunit_exec_fast_alu_result_to_writeback_pipe_read_ack : out std_logic_vector(0 downto 0);
    iunit_exec_to_writeback_pipe_read_data: out std_logic_vector(125 downto 0);
    iunit_exec_to_writeback_pipe_read_req : in std_logic_vector(0 downto 0);
    iunit_exec_to_writeback_pipe_read_ack : out std_logic_vector(0 downto 0);
    iunit_register_file_read_access_response_pipe_write_data: in std_logic_vector(141 downto 0);
    iunit_register_file_read_access_response_pipe_write_req : in std_logic_vector(0 downto 0);
    iunit_register_file_read_access_response_pipe_write_ack : out std_logic_vector(0 downto 0);
    noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_read_data: out std_logic_vector(16 downto 0);
    noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_read_req : in std_logic_vector(0 downto 0);
    noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_read_ack : out std_logic_vector(0 downto 0);
    noblock_iunit_exec_bypass_signal_to_register_file_pipe_read_data: out std_logic_vector(82 downto 0);
    noblock_iunit_exec_bypass_signal_to_register_file_pipe_read_req : in std_logic_vector(0 downto 0);
    noblock_iunit_exec_bypass_signal_to_register_file_pipe_read_ack : out std_logic_vector(0 downto 0);
    noblock_iunit_exec_to_regfile_credit_return_pipe_read_data: out std_logic_vector(0 downto 0);
    noblock_iunit_exec_to_regfile_credit_return_pipe_read_req : in std_logic_vector(0 downto 0);
    noblock_iunit_exec_to_regfile_credit_return_pipe_read_ack : out std_logic_vector(0 downto 0);
    teu_idispatch_to_iunit_exec_pipe_write_data: in std_logic_vector(149 downto 0);
    teu_idispatch_to_iunit_exec_pipe_write_req : in std_logic_vector(0 downto 0);
    teu_idispatch_to_iunit_exec_pipe_write_ack : out std_logic_vector(0 downto 0);
    teu_iunit_to_stream_corrector_pipe_read_data: out std_logic_vector(89 downto 0);
    teu_iunit_to_stream_corrector_pipe_read_req : in std_logic_vector(0 downto 0);
    teu_iunit_to_stream_corrector_pipe_read_ack : out std_logic_vector(0 downto 0);
    teu_iunit_trap_to_fpunit_pipe_read_data: out std_logic_vector(12 downto 0);
    teu_iunit_trap_to_fpunit_pipe_read_req : in std_logic_vector(0 downto 0);
    teu_iunit_trap_to_fpunit_pipe_read_ack : out std_logic_vector(0 downto 0);
    teu_iunit_trap_to_loadstore_pipe_read_data: out std_logic_vector(0 downto 0);
    teu_iunit_trap_to_loadstore_pipe_read_req : in std_logic_vector(0 downto 0);
    teu_iunit_trap_to_loadstore_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture iu_exec_arch  of iu_exec is -- system-architecture 
  -- interface signals to connect to memory space memory_space_1
  -- declarations related to module alignDivisorToDividendRevised
  -- declarations related to module decode_alu_exec_control_word
  -- declarations related to module exec_cti_instruction
  -- declarations related to module exec_eval_icc
  -- declarations related to module exec_rett_instruction
  -- declarations related to module find_left_16
  -- declarations related to module find_left_32
  -- declarations related to module find_left_4
  -- declarations related to module find_left_8
  -- declarations related to module find_leftmost_64
  -- declarations related to module i32_add_sub
  -- declarations related to module i32_div
  component i32_div is -- 
    generic (tag_length : integer); 
    port ( -- 
      signed_div : in  std_logic_vector(0 downto 0);
      set_cc : in  std_logic_vector(0 downto 0);
      y_in : in  std_logic_vector(31 downto 0);
      dividend : in  std_logic_vector(31 downto 0);
      divisor : in  std_logic_vector(31 downto 0);
      result : out  std_logic_vector(31 downto 0);
      No : out  std_logic_vector(0 downto 0);
      Zo : out  std_logic_vector(0 downto 0);
      Vo : out  std_logic_vector(0 downto 0);
      Co : out  std_logic_vector(0 downto 0);
      u64_true_divide_revised_call_reqs : out  std_logic_vector(0 downto 0);
      u64_true_divide_revised_call_acks : in   std_logic_vector(0 downto 0);
      u64_true_divide_revised_call_data : out  std_logic_vector(95 downto 0);
      u64_true_divide_revised_call_tag  :  out  std_logic_vector(0 downto 0);
      u64_true_divide_revised_return_reqs : out  std_logic_vector(0 downto 0);
      u64_true_divide_revised_return_acks : in   std_logic_vector(0 downto 0);
      u64_true_divide_revised_return_data : in   std_logic_vector(63 downto 0);
      u64_true_divide_revised_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module i32_div
  signal i32_div_signed_div :  std_logic_vector(0 downto 0);
  signal i32_div_set_cc :  std_logic_vector(0 downto 0);
  signal i32_div_y_in :  std_logic_vector(31 downto 0);
  signal i32_div_dividend :  std_logic_vector(31 downto 0);
  signal i32_div_divisor :  std_logic_vector(31 downto 0);
  signal i32_div_result :  std_logic_vector(31 downto 0);
  signal i32_div_No :  std_logic_vector(0 downto 0);
  signal i32_div_Zo :  std_logic_vector(0 downto 0);
  signal i32_div_Vo :  std_logic_vector(0 downto 0);
  signal i32_div_Co :  std_logic_vector(0 downto 0);
  signal i32_div_in_args    : std_logic_vector(97 downto 0);
  signal i32_div_out_args   : std_logic_vector(35 downto 0);
  signal i32_div_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal i32_div_tag_out   : std_logic_vector(1 downto 0);
  signal i32_div_start_req : std_logic;
  signal i32_div_start_ack : std_logic;
  signal i32_div_fin_req   : std_logic;
  signal i32_div_fin_ack : std_logic;
  -- caller side aggregated signals for module i32_div
  signal i32_div_call_reqs: std_logic_vector(0 downto 0);
  signal i32_div_call_acks: std_logic_vector(0 downto 0);
  signal i32_div_return_reqs: std_logic_vector(0 downto 0);
  signal i32_div_return_acks: std_logic_vector(0 downto 0);
  signal i32_div_call_data: std_logic_vector(97 downto 0);
  signal i32_div_call_tag: std_logic_vector(0 downto 0);
  signal i32_div_return_data: std_logic_vector(35 downto 0);
  signal i32_div_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module i32_mul_calculate_sign_correction
  -- declarations related to module i32_mulscc
  -- declarations related to module i32_shift
  -- declarations related to module i32_sll
  -- declarations related to module i32_srl
  -- declarations related to module increment_16
  -- declarations related to module increment_32
  -- declarations related to module increment_64
  -- declarations related to module increment_8
  -- declarations related to module iu_exec_daemon
  component iu_exec_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      iunit_register_file_read_access_response_pipe_read_req : out  std_logic_vector(0 downto 0);
      iunit_register_file_read_access_response_pipe_read_ack : in   std_logic_vector(0 downto 0);
      iunit_register_file_read_access_response_pipe_read_data : in   std_logic_vector(141 downto 0);
      teu_idispatch_to_iunit_exec_pipe_read_req : out  std_logic_vector(0 downto 0);
      teu_idispatch_to_iunit_exec_pipe_read_ack : in   std_logic_vector(0 downto 0);
      teu_idispatch_to_iunit_exec_pipe_read_data : in   std_logic_vector(149 downto 0);
      noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_data : out  std_logic_vector(16 downto 0);
      noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_data : out  std_logic_vector(82 downto 0);
      noblock_iunit_exec_to_regfile_credit_return_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_iunit_exec_to_regfile_credit_return_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_iunit_exec_to_regfile_credit_return_pipe_write_data : out  std_logic_vector(0 downto 0);
      iunit_exec_fast_alu_result_to_writeback_pipe_write_req : out  std_logic_vector(0 downto 0);
      iunit_exec_fast_alu_result_to_writeback_pipe_write_ack : in   std_logic_vector(0 downto 0);
      iunit_exec_fast_alu_result_to_writeback_pipe_write_data : out  std_logic_vector(108 downto 0);
      iunit_exec_to_writeback_pipe_write_req : out  std_logic_vector(0 downto 0);
      iunit_exec_to_writeback_pipe_write_ack : in   std_logic_vector(0 downto 0);
      iunit_exec_to_writeback_pipe_write_data : out  std_logic_vector(125 downto 0);
      teu_iunit_to_stream_corrector_pipe_write_req : out  std_logic_vector(0 downto 0);
      teu_iunit_to_stream_corrector_pipe_write_ack : in   std_logic_vector(0 downto 0);
      teu_iunit_to_stream_corrector_pipe_write_data : out  std_logic_vector(89 downto 0);
      teu_iunit_trap_to_fpunit_pipe_write_req : out  std_logic_vector(0 downto 0);
      teu_iunit_trap_to_fpunit_pipe_write_ack : in   std_logic_vector(0 downto 0);
      teu_iunit_trap_to_fpunit_pipe_write_data : out  std_logic_vector(12 downto 0);
      teu_iunit_trap_to_loadstore_pipe_write_req : out  std_logic_vector(0 downto 0);
      teu_iunit_trap_to_loadstore_pipe_write_ack : in   std_logic_vector(0 downto 0);
      teu_iunit_trap_to_loadstore_pipe_write_data : out  std_logic_vector(0 downto 0);
      i32_div_call_reqs : out  std_logic_vector(0 downto 0);
      i32_div_call_acks : in   std_logic_vector(0 downto 0);
      i32_div_call_data : out  std_logic_vector(97 downto 0);
      i32_div_call_tag  :  out  std_logic_vector(0 downto 0);
      i32_div_return_reqs : out  std_logic_vector(0 downto 0);
      i32_div_return_acks : in   std_logic_vector(0 downto 0);
      i32_div_return_data : in   std_logic_vector(35 downto 0);
      i32_div_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module iu_exec_daemon
  signal iu_exec_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal iu_exec_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal iu_exec_daemon_start_req : std_logic;
  signal iu_exec_daemon_start_ack : std_logic;
  signal iu_exec_daemon_fin_req   : std_logic;
  signal iu_exec_daemon_fin_ack : std_logic;
  -- declarations related to module iu_umul32
  -- declarations related to module restore_window_trap
  -- declarations related to module save_window_trap
  -- declarations related to module twos_complement_32
  -- declarations related to module twos_complement_64
  -- declarations related to module u32_sll
  -- declarations related to module u64_sll
  -- declarations related to module u64_true_divide_revised
  component u64_true_divide_revised is -- 
    generic (tag_length : integer); 
    port ( -- 
      udividend : in  std_logic_vector(63 downto 0);
      udivisor : in  std_logic_vector(31 downto 0);
      quotient : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module u64_true_divide_revised
  signal u64_true_divide_revised_udividend :  std_logic_vector(63 downto 0);
  signal u64_true_divide_revised_udivisor :  std_logic_vector(31 downto 0);
  signal u64_true_divide_revised_quotient :  std_logic_vector(63 downto 0);
  signal u64_true_divide_revised_in_args    : std_logic_vector(95 downto 0);
  signal u64_true_divide_revised_out_args   : std_logic_vector(63 downto 0);
  signal u64_true_divide_revised_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal u64_true_divide_revised_tag_out   : std_logic_vector(1 downto 0);
  signal u64_true_divide_revised_start_req : std_logic;
  signal u64_true_divide_revised_start_ack : std_logic;
  signal u64_true_divide_revised_fin_req   : std_logic;
  signal u64_true_divide_revised_fin_ack : std_logic;
  -- caller side aggregated signals for module u64_true_divide_revised
  signal u64_true_divide_revised_call_reqs: std_logic_vector(0 downto 0);
  signal u64_true_divide_revised_call_acks: std_logic_vector(0 downto 0);
  signal u64_true_divide_revised_return_reqs: std_logic_vector(0 downto 0);
  signal u64_true_divide_revised_return_acks: std_logic_vector(0 downto 0);
  signal u64_true_divide_revised_call_data: std_logic_vector(95 downto 0);
  signal u64_true_divide_revised_call_tag: std_logic_vector(0 downto 0);
  signal u64_true_divide_revised_return_data: std_logic_vector(63 downto 0);
  signal u64_true_divide_revised_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module u64_true_divide_revised_core
  -- declarations related to module u_cmp_32
  -- declarations related to module u_cmp_34
  -- declarations related to module u_set_index_64
  -- aggregate signals for write to pipe iunit_exec_fast_alu_result_to_writeback
  signal iunit_exec_fast_alu_result_to_writeback_pipe_write_data: std_logic_vector(108 downto 0);
  signal iunit_exec_fast_alu_result_to_writeback_pipe_write_req: std_logic_vector(0 downto 0);
  signal iunit_exec_fast_alu_result_to_writeback_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe iunit_exec_to_writeback
  signal iunit_exec_to_writeback_pipe_write_data: std_logic_vector(125 downto 0);
  signal iunit_exec_to_writeback_pipe_write_req: std_logic_vector(0 downto 0);
  signal iunit_exec_to_writeback_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe iunit_register_file_read_access_response
  signal iunit_register_file_read_access_response_pipe_read_data: std_logic_vector(141 downto 0);
  signal iunit_register_file_read_access_response_pipe_read_req: std_logic_vector(0 downto 0);
  signal iunit_register_file_read_access_response_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_iunit_exec_bypass_cc_signal_to_register_file
  signal noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_data: std_logic_vector(16 downto 0);
  signal noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_iunit_exec_bypass_signal_to_register_file
  signal noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_data: std_logic_vector(82 downto 0);
  signal noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_iunit_exec_to_regfile_credit_return
  signal noblock_iunit_exec_to_regfile_credit_return_pipe_write_data: std_logic_vector(0 downto 0);
  signal noblock_iunit_exec_to_regfile_credit_return_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_iunit_exec_to_regfile_credit_return_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe teu_idispatch_to_iunit_exec
  signal teu_idispatch_to_iunit_exec_pipe_read_data: std_logic_vector(149 downto 0);
  signal teu_idispatch_to_iunit_exec_pipe_read_req: std_logic_vector(0 downto 0);
  signal teu_idispatch_to_iunit_exec_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe teu_iunit_to_stream_corrector
  signal teu_iunit_to_stream_corrector_pipe_write_data: std_logic_vector(89 downto 0);
  signal teu_iunit_to_stream_corrector_pipe_write_req: std_logic_vector(0 downto 0);
  signal teu_iunit_to_stream_corrector_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe teu_iunit_trap_to_fpunit
  signal teu_iunit_trap_to_fpunit_pipe_write_data: std_logic_vector(12 downto 0);
  signal teu_iunit_trap_to_fpunit_pipe_write_req: std_logic_vector(0 downto 0);
  signal teu_iunit_trap_to_fpunit_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe teu_iunit_trap_to_loadstore
  signal teu_iunit_trap_to_loadstore_pipe_write_data: std_logic_vector(0 downto 0);
  signal teu_iunit_trap_to_loadstore_pipe_write_req: std_logic_vector(0 downto 0);
  signal teu_iunit_trap_to_loadstore_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module i32_div
  i32_div_signed_div <= i32_div_in_args(97 downto 97);
  i32_div_set_cc <= i32_div_in_args(96 downto 96);
  i32_div_y_in <= i32_div_in_args(95 downto 64);
  i32_div_dividend <= i32_div_in_args(63 downto 32);
  i32_div_divisor <= i32_div_in_args(31 downto 0);
  i32_div_out_args <= i32_div_result & i32_div_No & i32_div_Zo & i32_div_Vo & i32_div_Co ;
  -- call arbiter for module i32_div
  i32_div_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 98,
      return_data_width => 36,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => i32_div_call_reqs,
      call_acks => i32_div_call_acks,
      return_reqs => i32_div_return_reqs,
      return_acks => i32_div_return_acks,
      call_data  => i32_div_call_data,
      call_tag  => i32_div_call_tag,
      return_tag  => i32_div_return_tag,
      call_mtag => i32_div_tag_in,
      return_mtag => i32_div_tag_out,
      return_data =>i32_div_return_data,
      call_mreq => i32_div_start_req,
      call_mack => i32_div_start_ack,
      return_mreq => i32_div_fin_req,
      return_mack => i32_div_fin_ack,
      call_mdata => i32_div_in_args,
      return_mdata => i32_div_out_args,
      clk => clk, 
      reset => reset --
    ); --
  i32_div_instance:i32_div-- 
    generic map(tag_length => 2)
    port map(-- 
      signed_div => i32_div_signed_div,
      set_cc => i32_div_set_cc,
      y_in => i32_div_y_in,
      dividend => i32_div_dividend,
      divisor => i32_div_divisor,
      result => i32_div_result,
      No => i32_div_No,
      Zo => i32_div_Zo,
      Vo => i32_div_Vo,
      Co => i32_div_Co,
      start_req => i32_div_start_req,
      start_ack => i32_div_start_ack,
      fin_req => i32_div_fin_req,
      fin_ack => i32_div_fin_ack,
      clk => clk,
      reset => reset,
      u64_true_divide_revised_call_reqs => u64_true_divide_revised_call_reqs(0 downto 0),
      u64_true_divide_revised_call_acks => u64_true_divide_revised_call_acks(0 downto 0),
      u64_true_divide_revised_call_data => u64_true_divide_revised_call_data(95 downto 0),
      u64_true_divide_revised_call_tag => u64_true_divide_revised_call_tag(0 downto 0),
      u64_true_divide_revised_return_reqs => u64_true_divide_revised_return_reqs(0 downto 0),
      u64_true_divide_revised_return_acks => u64_true_divide_revised_return_acks(0 downto 0),
      u64_true_divide_revised_return_data => u64_true_divide_revised_return_data(63 downto 0),
      u64_true_divide_revised_return_tag => u64_true_divide_revised_return_tag(0 downto 0),
      tag_in => i32_div_tag_in,
      tag_out => i32_div_tag_out-- 
    ); -- 
  -- module iu_exec_daemon
  iu_exec_daemon_instance:iu_exec_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => iu_exec_daemon_start_req,
      start_ack => iu_exec_daemon_start_ack,
      fin_req => iu_exec_daemon_fin_req,
      fin_ack => iu_exec_daemon_fin_ack,
      clk => clk,
      reset => reset,
      iunit_register_file_read_access_response_pipe_read_req => iunit_register_file_read_access_response_pipe_read_req(0 downto 0),
      iunit_register_file_read_access_response_pipe_read_ack => iunit_register_file_read_access_response_pipe_read_ack(0 downto 0),
      iunit_register_file_read_access_response_pipe_read_data => iunit_register_file_read_access_response_pipe_read_data(141 downto 0),
      teu_idispatch_to_iunit_exec_pipe_read_req => teu_idispatch_to_iunit_exec_pipe_read_req(0 downto 0),
      teu_idispatch_to_iunit_exec_pipe_read_ack => teu_idispatch_to_iunit_exec_pipe_read_ack(0 downto 0),
      teu_idispatch_to_iunit_exec_pipe_read_data => teu_idispatch_to_iunit_exec_pipe_read_data(149 downto 0),
      noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_req => noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_req(0 downto 0),
      noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_ack => noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_ack(0 downto 0),
      noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_data => noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_data(16 downto 0),
      noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_req => noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_req(0 downto 0),
      noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_ack => noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_ack(0 downto 0),
      noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_data => noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_data(82 downto 0),
      noblock_iunit_exec_to_regfile_credit_return_pipe_write_req => noblock_iunit_exec_to_regfile_credit_return_pipe_write_req(0 downto 0),
      noblock_iunit_exec_to_regfile_credit_return_pipe_write_ack => noblock_iunit_exec_to_regfile_credit_return_pipe_write_ack(0 downto 0),
      noblock_iunit_exec_to_regfile_credit_return_pipe_write_data => noblock_iunit_exec_to_regfile_credit_return_pipe_write_data(0 downto 0),
      iunit_exec_fast_alu_result_to_writeback_pipe_write_req => iunit_exec_fast_alu_result_to_writeback_pipe_write_req(0 downto 0),
      iunit_exec_fast_alu_result_to_writeback_pipe_write_ack => iunit_exec_fast_alu_result_to_writeback_pipe_write_ack(0 downto 0),
      iunit_exec_fast_alu_result_to_writeback_pipe_write_data => iunit_exec_fast_alu_result_to_writeback_pipe_write_data(108 downto 0),
      iunit_exec_to_writeback_pipe_write_req => iunit_exec_to_writeback_pipe_write_req(0 downto 0),
      iunit_exec_to_writeback_pipe_write_ack => iunit_exec_to_writeback_pipe_write_ack(0 downto 0),
      iunit_exec_to_writeback_pipe_write_data => iunit_exec_to_writeback_pipe_write_data(125 downto 0),
      teu_iunit_to_stream_corrector_pipe_write_req => teu_iunit_to_stream_corrector_pipe_write_req(0 downto 0),
      teu_iunit_to_stream_corrector_pipe_write_ack => teu_iunit_to_stream_corrector_pipe_write_ack(0 downto 0),
      teu_iunit_to_stream_corrector_pipe_write_data => teu_iunit_to_stream_corrector_pipe_write_data(89 downto 0),
      teu_iunit_trap_to_fpunit_pipe_write_req => teu_iunit_trap_to_fpunit_pipe_write_req(0 downto 0),
      teu_iunit_trap_to_fpunit_pipe_write_ack => teu_iunit_trap_to_fpunit_pipe_write_ack(0 downto 0),
      teu_iunit_trap_to_fpunit_pipe_write_data => teu_iunit_trap_to_fpunit_pipe_write_data(12 downto 0),
      teu_iunit_trap_to_loadstore_pipe_write_req => teu_iunit_trap_to_loadstore_pipe_write_req(0 downto 0),
      teu_iunit_trap_to_loadstore_pipe_write_ack => teu_iunit_trap_to_loadstore_pipe_write_ack(0 downto 0),
      teu_iunit_trap_to_loadstore_pipe_write_data => teu_iunit_trap_to_loadstore_pipe_write_data(0 downto 0),
      i32_div_call_reqs => i32_div_call_reqs(0 downto 0),
      i32_div_call_acks => i32_div_call_acks(0 downto 0),
      i32_div_call_data => i32_div_call_data(97 downto 0),
      i32_div_call_tag => i32_div_call_tag(0 downto 0),
      i32_div_return_reqs => i32_div_return_reqs(0 downto 0),
      i32_div_return_acks => i32_div_return_acks(0 downto 0),
      i32_div_return_data => i32_div_return_data(35 downto 0),
      i32_div_return_tag => i32_div_return_tag(0 downto 0),
      tag_in => iu_exec_daemon_tag_in,
      tag_out => iu_exec_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  iu_exec_daemon_tag_in <= (others => '0');
  iu_exec_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => iu_exec_daemon_start_req, start_ack => iu_exec_daemon_start_ack,  fin_req => iu_exec_daemon_fin_req,  fin_ack => iu_exec_daemon_fin_ack);
  -- module u64_true_divide_revised
  u64_true_divide_revised_udividend <= u64_true_divide_revised_in_args(95 downto 32);
  u64_true_divide_revised_udivisor <= u64_true_divide_revised_in_args(31 downto 0);
  u64_true_divide_revised_out_args <= u64_true_divide_revised_quotient ;
  -- call arbiter for module u64_true_divide_revised
  u64_true_divide_revised_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 96,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => u64_true_divide_revised_call_reqs,
      call_acks => u64_true_divide_revised_call_acks,
      return_reqs => u64_true_divide_revised_return_reqs,
      return_acks => u64_true_divide_revised_return_acks,
      call_data  => u64_true_divide_revised_call_data,
      call_tag  => u64_true_divide_revised_call_tag,
      return_tag  => u64_true_divide_revised_return_tag,
      call_mtag => u64_true_divide_revised_tag_in,
      return_mtag => u64_true_divide_revised_tag_out,
      return_data =>u64_true_divide_revised_return_data,
      call_mreq => u64_true_divide_revised_start_req,
      call_mack => u64_true_divide_revised_start_ack,
      return_mreq => u64_true_divide_revised_fin_req,
      return_mack => u64_true_divide_revised_fin_ack,
      call_mdata => u64_true_divide_revised_in_args,
      return_mdata => u64_true_divide_revised_out_args,
      clk => clk, 
      reset => reset --
    ); --
  u64_true_divide_revised_instance:u64_true_divide_revised-- 
    generic map(tag_length => 2)
    port map(-- 
      udividend => u64_true_divide_revised_udividend,
      udivisor => u64_true_divide_revised_udivisor,
      quotient => u64_true_divide_revised_quotient,
      start_req => u64_true_divide_revised_start_req,
      start_ack => u64_true_divide_revised_start_ack,
      fin_req => u64_true_divide_revised_fin_req,
      fin_ack => u64_true_divide_revised_fin_ack,
      clk => clk,
      reset => reset,
      tag_in => u64_true_divide_revised_tag_in,
      tag_out => u64_true_divide_revised_tag_out-- 
    ); -- 
  iunit_exec_fast_alu_result_to_writeback_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe iunit_exec_fast_alu_result_to_writeback",
      num_reads => 1,
      num_writes => 1,
      data_width => 109,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => iunit_exec_fast_alu_result_to_writeback_pipe_read_req,
      read_ack => iunit_exec_fast_alu_result_to_writeback_pipe_read_ack,
      read_data => iunit_exec_fast_alu_result_to_writeback_pipe_read_data,
      write_req => iunit_exec_fast_alu_result_to_writeback_pipe_write_req,
      write_ack => iunit_exec_fast_alu_result_to_writeback_pipe_write_ack,
      write_data => iunit_exec_fast_alu_result_to_writeback_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  iunit_exec_to_writeback_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe iunit_exec_to_writeback",
      num_reads => 1,
      num_writes => 1,
      data_width => 126,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => iunit_exec_to_writeback_pipe_read_req,
      read_ack => iunit_exec_to_writeback_pipe_read_ack,
      read_data => iunit_exec_to_writeback_pipe_read_data,
      write_req => iunit_exec_to_writeback_pipe_write_req,
      write_ack => iunit_exec_to_writeback_pipe_write_ack,
      write_data => iunit_exec_to_writeback_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  iunit_register_file_read_access_response_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe iunit_register_file_read_access_response",
      num_reads => 1,
      num_writes => 1,
      data_width => 142,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => iunit_register_file_read_access_response_pipe_read_req,
      read_ack => iunit_register_file_read_access_response_pipe_read_ack,
      read_data => iunit_register_file_read_access_response_pipe_read_data,
      write_req => iunit_register_file_read_access_response_pipe_write_req,
      write_ack => iunit_register_file_read_access_response_pipe_write_ack,
      write_data => iunit_register_file_read_access_response_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_iunit_exec_bypass_cc_signal_to_register_file_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_iunit_exec_bypass_cc_signal_to_register_file",
      num_reads => 1,
      num_writes => 1,
      data_width => 17,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_read_req,
      read_ack => noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_read_ack,
      read_data => noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_read_data,
      write_req => noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_req,
      write_ack => noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_ack,
      write_data => noblock_iunit_exec_bypass_cc_signal_to_register_file_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_iunit_exec_bypass_signal_to_register_file_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_iunit_exec_bypass_signal_to_register_file",
      num_reads => 1,
      num_writes => 1,
      data_width => 83,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => noblock_iunit_exec_bypass_signal_to_register_file_pipe_read_req,
      read_ack => noblock_iunit_exec_bypass_signal_to_register_file_pipe_read_ack,
      read_data => noblock_iunit_exec_bypass_signal_to_register_file_pipe_read_data,
      write_req => noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_req,
      write_ack => noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_ack,
      write_data => noblock_iunit_exec_bypass_signal_to_register_file_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_iunit_exec_to_regfile_credit_return_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_iunit_exec_to_regfile_credit_return",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => noblock_iunit_exec_to_regfile_credit_return_pipe_read_req,
      read_ack => noblock_iunit_exec_to_regfile_credit_return_pipe_read_ack,
      read_data => noblock_iunit_exec_to_regfile_credit_return_pipe_read_data,
      write_req => noblock_iunit_exec_to_regfile_credit_return_pipe_write_req,
      write_ack => noblock_iunit_exec_to_regfile_credit_return_pipe_write_ack,
      write_data => noblock_iunit_exec_to_regfile_credit_return_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  teu_idispatch_to_iunit_exec_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe teu_idispatch_to_iunit_exec",
      num_reads => 1,
      num_writes => 1,
      data_width => 150,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => teu_idispatch_to_iunit_exec_pipe_read_req,
      read_ack => teu_idispatch_to_iunit_exec_pipe_read_ack,
      read_data => teu_idispatch_to_iunit_exec_pipe_read_data,
      write_req => teu_idispatch_to_iunit_exec_pipe_write_req,
      write_ack => teu_idispatch_to_iunit_exec_pipe_write_ack,
      write_data => teu_idispatch_to_iunit_exec_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  teu_iunit_to_stream_corrector_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe teu_iunit_to_stream_corrector",
      num_reads => 1,
      num_writes => 1,
      data_width => 90,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => teu_iunit_to_stream_corrector_pipe_read_req,
      read_ack => teu_iunit_to_stream_corrector_pipe_read_ack,
      read_data => teu_iunit_to_stream_corrector_pipe_read_data,
      write_req => teu_iunit_to_stream_corrector_pipe_write_req,
      write_ack => teu_iunit_to_stream_corrector_pipe_write_ack,
      write_data => teu_iunit_to_stream_corrector_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  teu_iunit_trap_to_fpunit_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe teu_iunit_trap_to_fpunit",
      num_reads => 1,
      num_writes => 1,
      data_width => 13,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => teu_iunit_trap_to_fpunit_pipe_read_req,
      read_ack => teu_iunit_trap_to_fpunit_pipe_read_ack,
      read_data => teu_iunit_trap_to_fpunit_pipe_read_data,
      write_req => teu_iunit_trap_to_fpunit_pipe_write_req,
      write_ack => teu_iunit_trap_to_fpunit_pipe_write_ack,
      write_data => teu_iunit_trap_to_fpunit_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  teu_iunit_trap_to_loadstore_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe teu_iunit_trap_to_loadstore",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => teu_iunit_trap_to_loadstore_pipe_read_req,
      read_ack => teu_iunit_trap_to_loadstore_pipe_read_ack,
      read_data => teu_iunit_trap_to_loadstore_pipe_read_data,
      write_req => teu_iunit_trap_to_loadstore_pipe_write_req,
      write_ack => teu_iunit_trap_to_loadstore_pipe_write_ack,
      write_data => teu_iunit_trap_to_loadstore_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  -- 
end iu_exec_arch;
